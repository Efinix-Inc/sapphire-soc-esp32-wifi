module top_soc (
output		    jtagCtrl_tdi,
input		    jtagCtrl_tdo,
output		    jtagCtrl_enable,
output		    jtagCtrl_capture,
output		    jtagCtrl_shift,
output		    jtagCtrl_update,
output		    jtagCtrl_reset,
input		    ut_jtagCtrl_tdi,
output		    ut_jtagCtrl_tdo,
input		    ut_jtagCtrl_enable,
input		    ut_jtagCtrl_capture,
input		    ut_jtagCtrl_shift,
input		    ut_jtagCtrl_update,
input		    ut_jtagCtrl_reset,
input		    io_cfuClk,
input		    io_cfuReset,
input		    cpu0_customInstruction_cmd_valid,
output		    cpu0_customInstruction_cmd_ready,
input [9:0]     cpu0_customInstruction_function_id,
input [31:0]    cpu0_customInstruction_inputs_0,
input [31:0]    cpu0_customInstruction_inputs_1,
output		    cpu0_customInstruction_rsp_valid,
input		    cpu0_customInstruction_rsp_ready,
output [31:0]   cpu0_customInstruction_outputs_0,
input		    cpu1_customInstruction_cmd_valid,
output		    cpu1_customInstruction_cmd_ready,
input [9:0]     cpu1_customInstruction_function_id,
input [31:0]    cpu1_customInstruction_inputs_0,
input [31:0]    cpu1_customInstruction_inputs_1,
output		    cpu1_customInstruction_rsp_valid,
input		    cpu1_customInstruction_rsp_ready,
output [31:0]   cpu1_customInstruction_outputs_0,
input		    cpu2_customInstruction_cmd_valid,
output		    cpu2_customInstruction_cmd_ready,
input [9:0]     cpu2_customInstruction_function_id,
input [31:0]    cpu2_customInstruction_inputs_0,
input [31:0]    cpu2_customInstruction_inputs_1,
output		    cpu2_customInstruction_rsp_valid,
input		    cpu2_customInstruction_rsp_ready,
output [31:0]   cpu2_customInstruction_outputs_0,
input		    cpu3_customInstruction_cmd_valid,
output		    cpu3_customInstruction_cmd_ready,
input [9:0]     cpu3_customInstruction_function_id,
input [31:0]    cpu3_customInstruction_inputs_0,
input [31:0]    cpu3_customInstruction_inputs_1,
output		    cpu3_customInstruction_rsp_valid,
input		    cpu3_customInstruction_rsp_ready,
output [31:0]   cpu3_customInstruction_outputs_0,
output		    io_ddrMasters_0_aw_valid,
input		    io_ddrMasters_0_aw_ready,
output [31:0]   io_ddrMasters_0_aw_payload_addr,
output [3:0]    io_ddrMasters_0_aw_payload_id,
output [3:0]    io_ddrMasters_0_aw_payload_region,
output [7:0]    io_ddrMasters_0_aw_payload_len,
output [2:0]    io_ddrMasters_0_aw_payload_size,
output [1:0]    io_ddrMasters_0_aw_payload_burst,
output		    io_ddrMasters_0_aw_payload_lock,
output [3:0]    io_ddrMasters_0_aw_payload_cache,
output [3:0]    io_ddrMasters_0_aw_payload_qos,
output [2:0]    io_ddrMasters_0_aw_payload_prot,
output		    io_ddrMasters_0_aw_payload_allStrb,
output		    io_ddrMasters_0_w_valid,
input		    io_ddrMasters_0_w_ready,
output [127:0]  io_ddrMasters_0_w_payload_data,
output [15:0]   io_ddrMasters_0_w_payload_strb,
output		    io_ddrMasters_0_w_payload_last,
input		    io_ddrMasters_0_b_valid,
output		    io_ddrMasters_0_b_ready,
input [3:0]     io_ddrMasters_0_b_payload_id,
input [1:0]     io_ddrMasters_0_b_payload_resp,
output		    io_ddrMasters_0_ar_valid,
input		    io_ddrMasters_0_ar_ready,
output [31:0]   io_ddrMasters_0_ar_payload_addr,
output [3:0]    io_ddrMasters_0_ar_payload_id,
output [3:0]    io_ddrMasters_0_ar_payload_region,
output [7:0]    io_ddrMasters_0_ar_payload_len,
output [2:0]    io_ddrMasters_0_ar_payload_size,
output [1:0]    io_ddrMasters_0_ar_payload_burst,
output		    io_ddrMasters_0_ar_payload_lock,
output [3:0]    io_ddrMasters_0_ar_payload_cache,
output [3:0]    io_ddrMasters_0_ar_payload_qos,
output [2:0]    io_ddrMasters_0_ar_payload_prot,
input		    io_ddrMasters_0_r_valid,
output		    io_ddrMasters_0_r_ready,
input [127:0]   io_ddrMasters_0_r_payload_data,
input [3:0]     io_ddrMasters_0_r_payload_id,
input [1:0]     io_ddrMasters_0_r_payload_resp,
input		    io_ddrMasters_0_r_payload_last,
input		    io_ddrMasters_0_clk,
input		    io_ddrMasters_0_reset,
output          io_ddrMasters_memCheck_pass,
output		    userInterruptA,
output		    userInterruptB,
output		    userInterruptC,
output		    userInterruptD,
output		    userInterruptE,
output		    userInterruptF,
output		    userInterruptH,
output		    userInterruptG,
output          userInterruptI,
output          userInterruptJ,
input [3:0]     system_gpio_0_io_read,
output [3:0]    system_gpio_0_io_write,
output [3:0]    system_gpio_0_io_writeEnable,
output		    system_uart_0_io_txd,
input		    system_uart_0_io_rxd,
output		    system_spi_0_io_sclk_write,
output		    system_spi_0_io_data_0_writeEnable,
input		    system_spi_0_io_data_0_read,
output		    system_spi_0_io_data_0_write,
output		    system_spi_0_io_data_1_writeEnable,
input		    system_spi_0_io_data_1_read,
output		    system_spi_0_io_data_1_write,
output		    system_spi_0_io_data_2_writeEnable,
input		    system_spi_0_io_data_2_read,
output		    system_spi_0_io_data_2_write,
output		    system_spi_0_io_data_3_writeEnable,
input		    system_spi_0_io_data_3_read,
output		    system_spi_0_io_data_3_write,
output [3:0]    system_spi_0_io_ss,
output		    system_i2c_0_io_sda_writeEnable,
output		    system_i2c_0_io_sda_write,
input		    system_i2c_0_io_sda_read,
output		    system_i2c_0_io_scl_writeEnable,
output		    system_i2c_0_io_scl_write,
input		    system_i2c_0_io_scl_read,
input [31:0]    axiA_awaddr,
input [7:0]	    axiA_awlen,
input [2:0]	    axiA_awsize,
input [1:0]	    axiA_awburst,
input		    axiA_awlock,
input [3:0]	    axiA_awcache,
input [2:0]	    axiA_awprot,
input [3:0]	    axiA_awqos,
input [3:0]	    axiA_awregion,
input		    axiA_awvalid,
output		    axiA_awready,
input [31:0]    axiA_wdata,
input [3:0]     axiA_wstrb,
input		    axiA_wvalid,
input		    axiA_wlast,
output		    axiA_wready,
output [1:0]    axiA_bresp,
output		    axiA_bvalid,
input		    axiA_bready,
input [31:0]    axiA_araddr,
input [7:0]	    axiA_arlen,
input [2:0]	    axiA_arsize,
input [1:0]	    axiA_arburst,
input		    axiA_arlock,
input [3:0]	    axiA_arcache,
input [2:0]	    axiA_arprot,
input [3:0]	    axiA_arqos,
input [3:0]	    axiA_arregion,
input		    axiA_arvalid,
output		    axiA_arready,
output [31:0]   axiA_rdata,
output [1:0]    axiA_rresp,
output		    axiA_rlast,
output		    axiA_rvalid,
input		    axiA_rready,
output          axiAInterrupt,
input           cfg_done,
output          cfg_start,
output          cfg_sel,
output          cfg_reset,
input		    io_peripheralClk,
input           io_peripheralReset,
output          io_asyncReset,
input           io_gpio_sw_n, 
input           pll_peripheral_locked,
input           pll_system_locked,
input           esp_ready_n,
input  [3:0]    qspi_d_IN,
output [3:0]    qspi_d_OUT,
output [3:0]    qspi_d_OE,
output          qspi_sclk,
output          qspi_ss
);
////////////////////////////////////////////////////////////////////////////
localparam PERI_FREQ = 200;
localparam AXIS_DEV  = 1;
localparam SLB  = 0;
////////////////////////////////////////////////////////////////////////////
//  Switch between peripheral and slb
wire [(AXIS_DEV*32)-1:0]    gAXIS_m_awaddr;
wire [(AXIS_DEV*8)-1:0]	    gAXIS_m_awlen;
wire [(AXIS_DEV*3)-1:0]	    gAXIS_m_awsize;
wire [(AXIS_DEV*2)-1:0]     gAXIS_m_awburst;
wire [(AXIS_DEV*2)-1:0]     gAXIS_m_awlock;
wire [(AXIS_DEV*4)-1:0]	    gAXIS_m_awcache;
wire [(AXIS_DEV*4)-1:0]	    gAXIS_m_awprot;
wire [(AXIS_DEV*4)-1:0]	    gAXIS_m_awqos;
wire [(AXIS_DEV*4)-1:0]	    gAXIS_m_awregion;
wire [AXIS_DEV-1:0]         gAXIS_m_awvalid;
wire [AXIS_DEV-1:0]         gAXIS_m_awready;
wire [(AXIS_DEV*32)-1:0]    gAXIS_m_wdata;
wire [(AXIS_DEV*4)-1:0]     gAXIS_m_wstrb;
wire [AXIS_DEV-1:0]         gAXIS_m_wvalid;
wire [AXIS_DEV-1:0]         gAXIS_m_wlast;
wire [AXIS_DEV-1:0]         gAXIS_m_wready;
wire [(AXIS_DEV*2)-1:0]     gAXIS_m_bresp;
wire [AXIS_DEV-1:0]         gAXIS_m_bvalid;
wire [AXIS_DEV-1:0]         gAXIS_m_bready;
wire [(AXIS_DEV*32)-1:0]    gAXIS_m_araddr;
wire [(AXIS_DEV*8)-1:0]	    gAXIS_m_arlen;
wire [(AXIS_DEV*3)-1:0]	    gAXIS_m_arsize;
wire [(AXIS_DEV*2)-1:0]	    gAXIS_m_arburst;
wire [(AXIS_DEV*2)-1:0]     gAXIS_m_arlock;
wire [(AXIS_DEV*4)-1:0]	    gAXIS_m_arcache;
wire [(AXIS_DEV*4)-1:0]	    gAXIS_m_arprot;
wire [(AXIS_DEV*4)-1:0]	    gAXIS_m_arqos;
wire [(AXIS_DEV*4)-1:0]	    gAXIS_m_arregion;
wire [AXIS_DEV-1:0]         gAXIS_m_arvalid;
wire [AXIS_DEV-1:0]         gAXIS_m_arready;
wire [(AXIS_DEV*32)-1:0]    gAXIS_m_rdata;
wire [(AXIS_DEV*2)-1:0]     gAXIS_m_rresp;
wire [AXIS_DEV-1:0]         gAXIS_m_rlast;
wire [AXIS_DEV-1:0]         gAXIS_m_rvalid;
wire [AXIS_DEV-1:0]         gAXIS_m_rready;

//reset
wire                        io_asyncReset_soc;
wire                        watchdog_reset;

gAXIS_1to3_switch u_AXIS_1to3_switch
(
    .rst_n              ( ~io_peripheralReset ),
    .clk                ( io_peripheralClk ),
    .m_axi_awvalid      ( gAXIS_m_awvalid ),
    .m_axi_awready      ( gAXIS_m_awready ),
    .m_axi_awid         ( ),
    .m_axi_awaddr       ( gAXIS_m_awaddr ),
    .m_axi_awburst      ( gAXIS_m_awburst ),
    .m_axi_awlen        ( gAXIS_m_awlen ),
    .m_axi_awsize       ( gAXIS_m_awsize ),
    .m_axi_awcache      ( gAXIS_m_awcache ),
    .m_axi_awqos        ( gAXIS_m_awqos ),
    .m_axi_awprot       ( gAXIS_m_awprot ),
    .m_axi_awuser       ( ),
    .m_axi_awlock       ( gAXIS_m_awlock ),
    .m_axi_awregion     ( gAXIS_m_awregion ),
    .m_axi_wvalid       ( gAXIS_m_wvalid ),
    .m_axi_wready       ( gAXIS_m_wready ),
    .m_axi_wdata        ( gAXIS_m_wdata ),
    .m_axi_wstrb        ( gAXIS_m_wstrb ),
    .m_axi_wlast        ( gAXIS_m_wlast ),
    .m_axi_wuser        ( ),
    .m_axi_bready       ( gAXIS_m_bready ),
    .m_axi_bvalid       ( gAXIS_m_bvalid ),
    .m_axi_bresp        ( gAXIS_m_bresp ),
    .m_axi_buser        ( {AXIS_DEV{3'h0}} ),
    .m_axi_bid          ( {AXIS_DEV{8'h0}} ),
    .m_axi_arvalid      ( gAXIS_m_arvalid ),
    .m_axi_arready      ( gAXIS_m_arready ),
    .m_axi_arid         ( ),
    .m_axi_araddr       ( gAXIS_m_araddr ),
    .m_axi_arburst      ( gAXIS_m_arburst ),
    .m_axi_arlen        ( gAXIS_m_arlen ),
    .m_axi_arsize       ( gAXIS_m_arsize ),
    .m_axi_arlock       ( gAXIS_m_arlock ),
    .m_axi_arprot       ( gAXIS_m_arprot ),
    .m_axi_arcache      ( gAXIS_m_arcache ),
    .m_axi_arqos        ( gAXIS_m_arqos ),
    .m_axi_aruser       ( ),
    .m_axi_arregion     ( gAXIS_m_arregion ),
    .m_axi_ruser        ( {AXIS_DEV{3'h0}}),
    .m_axi_rvalid       ( gAXIS_m_rvalid ),
    .m_axi_rready       ( gAXIS_m_rready ),
    .m_axi_rid          ( {AXIS_DEV{8'h0}}),
    .m_axi_rdata        ( gAXIS_m_rdata ),
    .m_axi_rresp        ( gAXIS_m_rresp ),
    .m_axi_rlast        ( gAXIS_m_rlast ),
    .s_axi_awvalid      ( axiA_awvalid ),
    .s_axi_awready      ( axiA_awready ),
    .s_axi_awaddr       ( {7'h00, axiA_awaddr[24:0]} ),
    .s_axi_awid         ( 8'h00 ),
    .s_axi_awburst      ( axiA_awburst ),
    .s_axi_awlen        ( axiA_awlen ),
    .s_axi_awsize       ( axiA_awsize ),
    .s_axi_awprot       ( {1'b0, axiA_awprot} ),
    .s_axi_awlock       ( {1'b0, axiA_awlock} ),
    .s_axi_awcache      ( axiA_awcache ),
    .s_axi_awqos        ( axiA_awqos ),
    .s_axi_awuser       ( 3'h0 ),
    .s_axi_wvalid       ( axiA_wvalid ),
    .s_axi_wready       ( axiA_wready ),
    .s_axi_wid          ( 8'h00 ),
    .s_axi_wdata        ( axiA_wdata ),
    .s_axi_wlast        ( axiA_wlast ),
    .s_axi_wstrb        ( axiA_wstrb ),
    .s_axi_wuser        ( 3'h0 ),
    .s_axi_bvalid       ( axiA_bvalid ),
    .s_axi_bready       ( axiA_bready ),
    .s_axi_bresp        ( axiA_bresp ),
    .s_axi_bid          ( ),
    .s_axi_buser        ( ),
    .s_axi_arvalid      ( axiA_arvalid ),
    .s_axi_arready      ( axiA_arready ),
    .s_axi_araddr       ( {7'h00, axiA_araddr[24:0]} ),
    .s_axi_arid         ( 8'h00 ),
    .s_axi_arburst      ( axiA_arburst ),
    .s_axi_arlen        ( axiA_arlen ),
    .s_axi_arsize       ( axiA_arsize ),
    .s_axi_arprot       ( { 1'b0, axiA_arprot} ),
    .s_axi_arlock       ( { 1'b0, axiA_arlock} ),
    .s_axi_arcache      ( axiA_arcache ),
    .s_axi_arqos        ( axiA_arqos ),
    .s_axi_aruser       ( 3'h0 ),
    .s_axi_rready       ( axiA_rready ),
    .s_axi_rvalid       ( axiA_rvalid ),
    .s_axi_rdata        ( axiA_rdata ),
    .s_axi_rresp        ( axiA_rresp ),
    .s_axi_rlast        ( axiA_rlast ),
    .s_axi_rid          ( ),
    .s_axi_ruser        ( )
);

//spi dma
  
wire [7:0]    apb_spi_dma_PADDR;
wire [0:0]    apb_spi_dma_PSEL;
wire          apb_spi_dma_PENABLE;
wire          apb_spi_dma_PREADY;
wire          apb_spi_dma_PWRITE;
wire [31:0]   apb_spi_dma_PWDATA;
wire [31:0]   apb_spi_dma_PRDATA;

assign userInterruptJ = ~esp_ready_n;
Apb3SpiXdrMasterDmaCtrl spi_dma_inst(
.apb_PADDR              (apb_spi_dma_PADDR  ), 
.apb_PSEL               (apb_spi_dma_PSEL   ), 
.apb_PENABLE            (apb_spi_dma_PENABLE), 
.apb_PREADY             (apb_spi_dma_PREADY ), 
.apb_PWRITE             (apb_spi_dma_PWRITE ), 
.apb_PWDATA             (apb_spi_dma_PWDATA ), 
.apb_PRDATA             (apb_spi_dma_PRDATA ),

.axim_awvalid           (io_ddrMasters_0_aw_valid         ), 
.axim_awready           (io_ddrMasters_0_aw_ready         ), 
.axim_awaddr            (io_ddrMasters_0_aw_payload_addr  ), 
.axim_awid              (io_ddrMasters_0_aw_payload_id    ), 
.axim_awregion          (io_ddrMasters_0_aw_payload_region), 
.axim_awlen             (io_ddrMasters_0_aw_payload_len   ), 
.axim_awsize            (io_ddrMasters_0_aw_payload_size  ), 
.axim_awburst           (io_ddrMasters_0_aw_payload_burst ), 
.axim_awlock            (io_ddrMasters_0_aw_payload_lock  ), 
.axim_awcache           (io_ddrMasters_0_aw_payload_cache ), 
.axim_awqos             (io_ddrMasters_0_aw_payload_qos   ), 
.axim_awprot            (io_ddrMasters_0_aw_payload_prot  ), 
.axim_wvalid            (io_ddrMasters_0_w_valid          ), 
.axim_wready            (io_ddrMasters_0_w_ready          ), 
.axim_wdata             (io_ddrMasters_0_w_payload_data   ), 
.axim_wstrb             (io_ddrMasters_0_w_payload_strb   ), 
.axim_wlast             (io_ddrMasters_0_w_payload_last   ), 
.axim_bvalid            (io_ddrMasters_0_b_valid          ), 
.axim_bready            (io_ddrMasters_0_b_ready          ), 
.axim_bid               (io_ddrMasters_0_b_payload_id     ), 
.axim_bresp             (io_ddrMasters_0_b_payload_resp   ), 
.axim_arvalid           (io_ddrMasters_0_ar_valid         ), 
.axim_arready           (io_ddrMasters_0_ar_ready         ), 
.axim_araddr            (io_ddrMasters_0_ar_payload_addr  ), 
.axim_arid              (io_ddrMasters_0_ar_payload_id    ), 
.axim_arregion          (io_ddrMasters_0_ar_payload_region), 
.axim_arlen             (io_ddrMasters_0_ar_payload_len   ), 
.axim_arsize            (io_ddrMasters_0_ar_payload_size  ), 
.axim_arburst           (io_ddrMasters_0_ar_payload_burst ), 
.axim_arlock            (io_ddrMasters_0_ar_payload_lock  ), 
.axim_arcache           (io_ddrMasters_0_ar_payload_cache ), 
.axim_arqos             (io_ddrMasters_0_ar_payload_qos   ), 
.axim_arprot            (io_ddrMasters_0_ar_payload_prot  ), 
.axim_rvalid            (io_ddrMasters_0_r_valid          ), 
.axim_rready            (io_ddrMasters_0_r_ready          ), 
.axim_rdata             (io_ddrMasters_0_r_payload_data   ), 
.axim_rid               (io_ddrMasters_0_r_payload_id     ), 
.axim_rresp             (io_ddrMasters_0_r_payload_resp   ), 
.axim_rlast             (io_ddrMasters_0_r_payload_last   ),


.spi_sclk_write         ( qspi_sclk         ),
.spi_data_0_writeEnable ( qspi_d_OE[0]      ),
.spi_data_0_read        ( qspi_d_IN[0]      ),
.spi_data_0_write       ( qspi_d_OUT[0]     ),
.spi_data_1_writeEnable ( qspi_d_OE[1]      ),
.spi_data_1_read        ( qspi_d_IN[1]      ),
.spi_data_1_write       ( qspi_d_OUT[1]     ),
.spi_data_2_writeEnable ( qspi_d_OE[2]      ),
.spi_data_2_read        ( qspi_d_IN[2]      ),
.spi_data_2_write       ( qspi_d_OUT[2]     ),
.spi_data_3_writeEnable ( qspi_d_OE[3]      ),
.spi_data_3_read        ( qspi_d_IN[3]      ),
.spi_data_3_write       ( qspi_d_OUT[3]     ),
.spi_ss                 ( qspi_ss           ),


.intr                   ( intr              ),
.ctrl_clk               ( io_peripheralClk  ), 
.ctrl_reset             ( io_peripheralReset),
.clk                    ( io_ddrMasters_0_clk), 
.reset                  ( io_ddrMasters_0_reset)
);


assign io_asyncReset = io_asyncReset_soc | watchdog_reset; 

//axi4 bridge to various I/O
EfxSapphireHpSoc_slb u_top_peripherals(
.io_apbSlave_0_PADDR                    ( dma_apb3_paddr    ),
.io_apbSlave_0_PENABLE                  ( dma_apb3_penable  ),
.io_apbSlave_0_PRDATA                   ( dma_apb3_prdata   ),
.io_apbSlave_0_PREADY                   ( dma_apb3_pready   ),
.io_apbSlave_0_PSEL                     ( dma_apb3_psel     ),
.io_apbSlave_0_PSLVERROR                ( dma_apb3_pslverror),
.io_apbSlave_0_PWDATA                   ( dma_apb3_pwdata   ),
.io_apbSlave_0_PWRITE                   ( dma_apb3_pwrite   ),

.io_apbSlave_1_PADDR                    ( apb_spi_dma_PADDR  ),
.io_apbSlave_1_PENABLE                  ( apb_spi_dma_PENABLE),
.io_apbSlave_1_PRDATA                   ( apb_spi_dma_PRDATA ),
.io_apbSlave_1_PREADY                   ( apb_spi_dma_PREADY ),
.io_apbSlave_1_PSEL                     ( apb_spi_dma_PSEL   ),
.io_apbSlave_1_PWDATA                   ( apb_spi_dma_PWDATA ),
.io_apbSlave_1_PWRITE                   ( apb_spi_dma_PWRITE ),

.system_uart_0_io_txd                   ( system_uart_0_io_txd ),
.system_uart_0_io_rxd                   ( system_uart_0_io_rxd ),
.system_i2c_0_io_sda_writeEnable        ( system_i2c_0_io_sda_writeEnable ),
.system_i2c_0_io_sda_write              ( system_i2c_0_io_sda_write ),
.system_i2c_0_io_sda_read               ( system_i2c_0_io_sda_read ),
.system_i2c_0_io_scl_writeEnable        ( system_i2c_0_io_scl_writeEnable ),
.system_i2c_0_io_scl_write              ( system_i2c_0_io_scl_write ),
.system_i2c_0_io_scl_read               ( system_i2c_0_io_scl_read ),
.jtagCtrl_tdi                           ( jtagCtrl_tdi ),
.jtagCtrl_tdo                           ( jtagCtrl_tdo ),
.jtagCtrl_enable                        ( jtagCtrl_enable ),
.jtagCtrl_capture                       ( jtagCtrl_capture ),
.jtagCtrl_shift                         ( jtagCtrl_shift ),
.jtagCtrl_update                        ( jtagCtrl_update ),
.jtagCtrl_reset                         ( jtagCtrl_reset ),
.ut_jtagCtrl_tdi                        ( ut_jtagCtrl_tdi ),
.ut_jtagCtrl_tdo                        ( ut_jtagCtrl_tdo ),
.ut_jtagCtrl_enable                     ( ut_jtagCtrl_enable ),
.ut_jtagCtrl_capture                    ( ut_jtagCtrl_capture ),
.ut_jtagCtrl_shift                      ( ut_jtagCtrl_shift ),
.ut_jtagCtrl_update                     ( ut_jtagCtrl_update ),
.ut_jtagCtrl_reset                      ( ut_jtagCtrl_reset ),
.system_gpio_0_io_read                  ( system_gpio_0_io_read ),
.system_gpio_0_io_write                 ( system_gpio_0_io_write ),
.system_gpio_0_io_writeEnable           ( system_gpio_0_io_writeEnable ),
.system_watchdog_hardPanic_reset        ( watchdog_reset ),
.userInterruptA                         ( userInterruptA ),
.userInterruptB                         ( userInterruptB ),
.userInterruptC                         ( userInterruptC ),
.userInterruptD                         ( userInterruptD ),
.userInterruptE                         ( userInterruptE ),
.userInterruptF                         ( userInterruptF ),
.axiA_awvalid                           ( gAXIS_m_awvalid[SLB*1 +: 1] ),
.axiA_awready                           ( gAXIS_m_awready[SLB*1 +: 1] ),
.axiA_awaddr                            ( gAXIS_m_awaddr[SLB*32 +: 32] ),
.axiA_awlen                             ( gAXIS_m_awlen[SLB*8 +: 8] ),
.axiA_awburst                           ( gAXIS_m_awburst[SLB*2 +: 2] ),
.axiA_awsize                            ( gAXIS_m_awsize[SLB*3 +: 3] ),
.axiA_awcache                           ( gAXIS_m_awcache[SLB*4 +: 4] ),
.axiA_awprot                            ( gAXIS_m_awprot[SLB*3 +: 3] ),
.axiA_wvalid                            ( gAXIS_m_wvalid[SLB*1 +: 1] ),
.axiA_wready                            ( gAXIS_m_wready[SLB*1 +: 1] ),
.axiA_wdata                             ( gAXIS_m_wdata[SLB*32 +: 32] ),
.axiA_wstrb                             ( gAXIS_m_wstrb[SLB*4 +: 4] ),
.axiA_wlast                             ( gAXIS_m_wlast[SLB*1 +: 1] ),
.axiA_bvalid                            ( gAXIS_m_bvalid[SLB*1 +: 1] ),
.axiA_bready                            ( gAXIS_m_bready[SLB*1 +: 1] ),
.axiA_bresp                             ( gAXIS_m_bresp[SLB*2 +: 2] ),
.axiA_arvalid                           ( gAXIS_m_arvalid[SLB*1 +: 1] ),
.axiA_arready                           ( gAXIS_m_arready[SLB*1 +: 1] ),
.axiA_araddr                            ( gAXIS_m_araddr[SLB*32 +: 32] ),
.axiA_arlen                             ( gAXIS_m_arlen[SLB*8 +: 8] ),
.axiA_arburst                           ( gAXIS_m_arburst[SLB*2 +: 2]),
.axiA_arsize                            ( gAXIS_m_arsize[SLB*3 +: 3] ),
.axiA_arcache                           ( gAXIS_m_arcache[SLB*4 +: 4] ),
.axiA_arprot                            ( gAXIS_m_arprot[SLB*3 +: 3] ),
.axiA_rvalid                            ( gAXIS_m_rvalid[SLB*1 +: 1] ),
.axiA_rready                            ( gAXIS_m_rready[SLB*1 +: 1] ),
.axiA_rdata                             ( gAXIS_m_rdata[SLB*32 +: 32] ),
.axiA_rresp                             ( gAXIS_m_rresp[SLB*2 +: 2] ),
.axiA_rlast                             ( gAXIS_m_rlast[SLB*1 +: 1] ),
.axiAInterrupt                          ( axiAInterrupt ),
.cfg_done                               ( cfg_done ),
.cfg_start                              ( cfg_start ),
.cfg_sel                                ( cfg_sel ),
.cfg_reset                              ( cfg_reset ),
.io_peripheralClk                       ( io_peripheralClk ),
.io_peripheralReset                     ( io_peripheralReset ),
.io_asyncReset                          ( io_asyncReset_soc ),
.io_gpio_sw_n                           ( io_gpio_sw_n ), 
.pll_peripheral_locked                  ( pll_peripheral_locked ),
.pll_system_locked                      ( pll_system_locked )
);

endmodule
