// Generator : SpinalHDL dev    git head : f89ba3384f643a2242caa7924e960fec1c38dd89
// Component : Apb3SpiXdrMasterDmaCtrl

`timescale 1ns/1ps

module Apb3SpiXdrMasterDmaCtrl (
  input  wire [7:0]    apb_PADDR,
  input  wire [0:0]    apb_PSEL,
  input  wire          apb_PENABLE,
  output wire          apb_PREADY,
  input  wire          apb_PWRITE,
  input  wire [31:0]   apb_PWDATA,
  output wire [31:0]   apb_PRDATA,
  output wire          axim_awvalid,
  input  wire          axim_awready,
  output wire [31:0]   axim_awaddr,
  output wire [3:0]    axim_awid,
  output wire [3:0]    axim_awregion,
  output wire [7:0]    axim_awlen,
  output wire [2:0]    axim_awsize,
  output wire [1:0]    axim_awburst,
  output wire [0:0]    axim_awlock,
  output wire [3:0]    axim_awcache,
  output wire [3:0]    axim_awqos,
  output wire [2:0]    axim_awprot,
  output wire          axim_wvalid,
  input  wire          axim_wready,
  output wire [127:0]  axim_wdata,
  output wire [15:0]   axim_wstrb,
  output wire          axim_wlast,
  input  wire          axim_bvalid,
  output wire          axim_bready,
  input  wire [3:0]    axim_bid,
  input  wire [1:0]    axim_bresp,
  output wire          axim_arvalid,
  input  wire          axim_arready,
  output wire [31:0]   axim_araddr,
  output wire [3:0]    axim_arid,
  output wire [3:0]    axim_arregion,
  output wire [7:0]    axim_arlen,
  output wire [2:0]    axim_arsize,
  output wire [1:0]    axim_arburst,
  output wire [0:0]    axim_arlock,
  output wire [3:0]    axim_arcache,
  output wire [3:0]    axim_arqos,
  output wire [2:0]    axim_arprot,
  input  wire          axim_rvalid,
  output wire          axim_rready,
  input  wire [127:0]  axim_rdata,
  input  wire [3:0]    axim_rid,
  input  wire [1:0]    axim_rresp,
  input  wire          axim_rlast,
  output wire [0:0]    spi_sclk_write,
  output wire          spi_data_0_writeEnable,
  input  wire [0:0]    spi_data_0_read,
  output wire [0:0]    spi_data_0_write,
  output wire          spi_data_1_writeEnable,
  input  wire [0:0]    spi_data_1_read,
  output wire [0:0]    spi_data_1_write,
  output wire          spi_data_2_writeEnable,
  input  wire [0:0]    spi_data_2_read,
  output wire [0:0]    spi_data_2_write,
  output wire          spi_data_3_writeEnable,
  input  wire [0:0]    spi_data_3_read,
  output wire [0:0]    spi_data_3_write,
  output wire [0:0]    spi_ss,
  output wire          intr,
  input  wire          clk,
  input  wire          reset,
  input  wire          ctrl_clk,
  input  wire          ctrl_reset
);

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="ipecrypt"
`pragma protect encrypt_agent_info="http://ipencrypter.com Version: 20.0.8"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"

`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_block
QH/ung1PaF1OP/281ww2ZORFP4dZTozvnpmefCDLeBtyHwGQZd8uY1tcXwSXiW47
35O0zeVBc3d3yp/L2VMFBotJ14zwhPvSUp1TMSAzI15WE/ntDlHYJol76DcWRWZI
3Lq+6/v9DUOk7aX6oJ0AHEX6A0+RRneyGWdVbLwz6tc=
`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_block
Bh7BRvr7QKWm859CBtS4eqWMsZUtbUyHI/l2L7xfZbFXWimI45co2+F9MTv929tc
sqT26LzGngZxzMfXOCvbk9d5BYBbWomATg2tJXg3zyyj+zxmsjHeVW9Aiq4zpSOo
ilJIgYllB36Go04vOCFR8weg7L25J4D6uY/dBNes2aq4U/uf1rI4jeOj4qJo/2oG
CGV1SnSdG4y/f7wbkxSwelPg9GZumMwxAcTPHWfUDZKWaXmuZJBxlaNRXUm9P2Rk
On06OqzH0lSrCXGzuCvc7hqnddXTlXjB4dylkzejsr9sJnrrWM8kYWTEu2C1NHwk
LyljWTkvQWLwOvfE5f4Ojw==
`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_block
qcr/ChYZdGO92dTpfRWK+CcnAYm4wbuxK8RI3AXkZA60fI+edVolfjKErj2VOaFb
QqBVQHja+rhvNoxl0763F27HG6l7ZLWMVjhNUzn3fMtJmTOYFm0T9Rr8D90/JTns
tEeyANidRaXoHgXjVZ38zIm/njTYTNWX5CUIn9K3FiM=
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_block
pvslIi9yRXBdddS1ieI4sWWcTTcDOu3hWhEWICNLFrIfctZgeo5IHdOXvzNGh5Fk
K95M57HhDcxzhNff4zCuPAbUmTZQcMZO1ZWbujkTkVEcMXJE4W7bqd/w5WWPSPkt
YMCAdgHB1y3KvQXCvk8cpweYCIFstjdYz5BCayEsu2/wATV7TxH3ZI6A79Z3zvul
ttRPmodOtTi/aQo8sD+JhUyApskp102oLMIoGLg1ua36No6GlAOa4qxfh4bfP5L4
zDSO7W/KlcVrUseNL+31e5aboiedqMnuk3XHMQvFwNna+1eYWkq6xoMxKF7GkQ1g
P8lNWrx7Sh/pCIBN0gft9g==
`pragma protect key_keyowner="Efinix Inc."
`pragma protect key_keyname="EFX_K01"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_block
RCGStWIatiPR9OkI2RF915+dyHIneWbqxdpInmOFbHUj5xgj7/5rrlBRSNdc5SQ3
EgjBM3/5FYFBVzhRh4spjzdpMPK8d3p3hJVIUreZYX7eUXOZEbyMyosIm6PmMLiV
Z8MRvGLP95HJK5zYtT0I9g1UFqiFDBBWtr33fDjhXNGZnDya1W+sT6LBV3w54c/8
hKnd421/NMcRjq2eikyE7/gSujQwQxPM1+05H1uLi6uFzAHFThzgJ64yDGPF/BN6
bDCk7tfWjtM0bthI8frSMcJXmzlRvMF6K8gNHfiWVeAKgTnjjOiOczC8YCRIFu9E
2dRPT3sGPwhWf4rD8ABcqw==
`pragma protect encoding=(enctype="base64", line_length=64, bytes=76608)
`pragma protect data_block
3CZUknNEISvonAMWpaHU4QYB3j9i6wGN6DhjYHb8XZI2tUz3lEELozzVsSZCu7YE
CoTvQcqv+/ms0nTaUW1xA6rPqM5dyUD1eUd0PSksH4LPZY4FsYAAMmYsxTIocLM1
WMwAxEEuZAzgopGmbBQ+cHIJkLwsTUMWtxa3tCImK1Dgj33Dfbi/rq4lpi2KIHT+
pgPWF4ybt8ZmxVlGBDUVB4Olvsr52KvuiQRa3lfRm9woZJzuXXVP/TRGHtH82sKc
Urs+u9bke6un2Gg/yjUt4/BpTVlboBjU+orjraUykfQLB7QhftTvhUHNwwoKnp7H
qTypN0eWhkLEdM7yXwJFmslevrJX9mmuHg6st9jQGIaXyZGmCBU4kNyG/qdMhAkY
sFMvuJ6L3xdO4iKK8KZAAimOcocgWsHjePYBE9gr10GNMKIhLOgvmHgVyJNUtIS4
4qSPZFVCbS9kmgj4Nw4lbmeXz0lG8AOG8rBOT/dl2ZJeDW8FhSq+pRQZbaheoEDn
ZjLcKpRUCkPEa1hKSjnlsIDKC9r1++5ZG1t6fRnRrQZvf7v1C8YVEo9JAcFB78g4
IUCLzB2ctwR/p6F3+9OF4tg/uymgr2Ub3RBX5ajjB6Dm/t0BfTy3aJsBcDhEoH20
ZtvCRYcMDGLh1fxXwu+nB8VDGmoLoSDYr5hDeg3FnYDxc3PM1yXNOcsfEhOzpYP9
C00pVBQg47dGdSC0FcCiN0gCg52GA5y+U73CPAzVbHwOQxfFa9W9WElPGJrLmu0v
hSZgdwsKl5OdoT7nJPUuNBx1FGcxKXTN06fILVc8jvDR7uFTIdKlIcPEFext1VY6
6sJn2GVL6CiTE+4PAwydvAYwdoWrcQaYtC1Y2WMi8+ldsPb/UEwfftWUXhEUacFc
x5QikMtFzwdyr05bdpqjS1rmb3oBc+eaNhJ82oEJBC7CShz2aNHa23IqGa9KVs2d
pEBXtgZc9iu/3l8BVI016JqCRkKFXzv7gPa4ROMRF3M8ZUj/vHpxVzOsKCx98VDL
Fnz7MsWYkInmZ5kY2j7pFHRidLBj5aXdNCrW2Ct6YyC2iIaNIVoCUPi0iaWWaVip
Qv7xeuzWhbVFDAhGP2cdpJi4XuGVjbtMvWwf0OELtVl+KYoZ5gwKGOemJxF48DRI
ZeqDqs2V1wMV4JpBAj21zgVxIAShoM1WEbNkZZ29aDXxcqOVELp7epHjapwr0ofn
k3Fwg7AMoN4uiEmNjcX0+fy7JMunYZzm+ImaevF68m56HUYs8A6NaVRHyMHR6tek
pOEyhnozY5OgLn5lyXz4fwct+CVyjUlUA2cY3wdLZFLDmGK/paB/HEtSEaPCnEep
5FvDa8SjtaQFloFkiQG+k4Geke3qX6HSl7rrAQ76IGCrnHin2p0bQhX+X0xWAhQo
yuvwkTI9BpXD/k4tYA2c6Nb02CSKql8fOcEGVFx4qghBidABubYaQL4164Hzp7JC
JWAPF4Y+sXfAX6DGb0iyYSdstWkMgvyt+/i+oK6SmxmeUE4z7KVB4bVMFyohEiV5
ZVp6fVWx0IbbTdL9268xB3XHDXX6bm+V7Tn6kzk89iVCWyKECsmSgm43PxkKhZxh
8diU5x+vKFlQHLcAw1ZLPWTAUjxADZaxNOjvijgr5Tbu4BnYYF1XrCU8uLb1H3T1
N8bxvR10Pyhr7PzKzOxlCeVIBqQqaTK749jXwNX8wZUyMMw2ticmnFpd+otFNFsd
/gJ8TJuMEmszxt/LuVx8OCePAuZg4/xnw+GDTj+SIAREurMUJ4Sv968wujVMcREH
PKnPF0emJCKTIIyViLqpBkZi5BI/GHxgSsf+gCTMKawaniotzzn+Q16co+mmmOO9
d/GUsmtkTrexRdizhesBaZ4dkTdaHnQpOWDUYcGAIkdw5hcsO7Og9IHLTSuY8cuh
2OydlSWHZF9/to3cGWUn+P1UucuyTEjCn5x4q/zI1istXgx4MPn30ZsiNUPbLWAh
fp4dFp64vyByt7qSI4YkHohquMPVmYc1WtZbkxi5RNuy1q6ys2kou1Pm4lQHf0jU
cWb7tr0d7z83AJhxv0QxmbFAYdLDk+JVGmcopbRfIq8QEz6Sau6kTwnTDIqBbBK8
EA+Q44pPNtc11UiNZjj2fvft+5dF81qhDF0OsMGsEbckLGTMYhuKv7130isGn6Iy
QfB7qtsfGgzvHWKrGmTMeNDdVDglDQOYsbaw/ZJLQYqAGJmsTxSkg59/tk0zU0Cz
aHZ/4h2miW6F/J05hpnrnlY/BAR3x7HoLaiHhw3maJaWqHfFz662bEF/c2Y0Zmy+
5pQRIw5B2UTwerLrKaUQDhRYzXv5CE0mjXIGbYLuONkA0YgdyO7YFiclNtbjD/AP
VOMLI+upaBuA+RkFCixJCJY0khVsJblJ4xjUOWey70qqEFgHLoxz26hhvVr3/Oyz
5WVigWoKmiShN9v1PTpQDdOtrKXGywzGPQ6UkS44MURId1F03qoi0BhD5gNxOH8F
TldRQ6A89siC2XTUv9VdlZ42rSeeuYKg9yO+w1If0vyjrYQjNXdem2o0rGopOQyP
EHMzfCCSOxu53+DADHkBGoXwWyUasF+9pzy3Idq3EMQTsPx/MtJC8B72EzkWb6xU
K5otwzEc+MwvXF3Jyk9pov2l5RVKdgY4SuU2/mactHOdKfzA9iDmZWBhcx1GZ4V3
fi4DC58NwYTnLDSsTqts3ae4pO/nA8Bdqj9ISKV8NpHmWe7EonZyB8g/XRXYyOs8
NHz4WNxXxDt4WwGXJsQ3j2Fra8r48pqEU+mxBYMPxjBYce3jiaDHQP34Htdl394z
XFCwHG/QVMkylI8x6Pr+JUlZP4WSq5GF9AtXTok8S191Xap88WKLI/GEwFHOgBR6
AkI/pd+XQJvPrDX5T6wtckImv4XNWgKtgpF/Nq/Lu/eUrPlELBrJ5PVefse/6CWO
T3+jzDAnWnSU8Rs4NNcBBTAN/Te9OkHF6knQnl7hQ7vxaUFX1MJjWsHXXZgR0O7Z
IZLB/Qpo2+Yj9TZk1SFZDNlWJuH+lL3HK89T8l+rQ3Sa1hCQKHpQcO2TVRYqNqzX
wqq9n0QFGlXCed1yEQ0Pwp5+3EzAbDhNommo3A95qUOekP6Cb5pnQPwAxyJND4Z/
dyXSQFCTP65EiOvVdVz5caS6xXq2W9yZfMbJjr37O5WTWpczY0v50hFA8/XazZe3
PXGspVZynUzn1tAHrd+6KPjDMOKzrk7vl8ulR5irM+gGotY0Y7sK2mhWYnPU/KL0
h8BIf7zbMMrO08C1Q5J3jeJc+4n9dDTAHtXmI2fwmWrVXLJhDGbtxDIzbxqIJIX/
eYWp3iC/Ho4e89DnMrM6nXEJOzg9i0+Bk54uaZ4Whg4RYwn8j5Zt3fBWosN5ERW2
zSXtU7IeiP5hdPeas3lK1OWrNWVj5VKbcFKREm4GtgJLtjdk9s9ECl9uGORvvyAh
4EkBnADRxX4+GC7z90W2tQZsYdP/ae0gN/nYtD3P08zyAdWDgGmNEuuCfEKmyxpx
n77M0z/AX1D5Iq9wHRY9GI7wn4mEs4aCMFiY9SrI00rIAvi2daMB2+0sEbpN0Poz
as8ot6Hvfd0uQM4Jp1wEptpJB2/WVukn0nK+aTbtIalIFsP88tn2mNpr8OCgdp/u
zSxTCI1mvVRZQGXKJxDdKoMykYG5zTAJUW1R89Lo7rBjA2bDCZx4dyR6rYaOK+Uz
5kN1wgcRYyDcRqjntJ73JcS4lZBnDU94LHTQMcl9lfGkc+n8fGmRuc/pUKPnp2wc
Y5ET0UfhAOu4QHB4BQi4L2RFqlLJxwtjayDE2mGpfuywjbd2OguXSV81OWjb1XEt
ecI/bDSnPv8sk+JDEhdI4sv21tagk5q4q9dQswqLnYeaGMWJ6/udA+xHF5K23HGP
3Ewpy6pkIAHu4+yxuIpMtSIHYJ0mt/GnUikrjcq13klklI3FduYdkKs9P4vtvWCY
SymajW+LNRQZpTgCcV6WXZMIxf3WsGzu1DlwPCilMfoYc6/9385t9e5/R5CwCkJn
K9eDTJT9+335F8cPhRHOC9b4dujhh8MHngdBq7mM2nwsLWKkFcKEzdmdf+o+Tebj
SRTg9WBY8Fh/9UsM0O2yEDWLOL5HaKvtY9MKwvGxpgsrqKSbs3NNKvtvRLxfw00N
106v1CffeVSD2MBBaeRr+azl4CjRWswCUxs/9VgjrkubIL1XUZ+wcVkzNjqSTYxP
J0cyUymdj4YlYtrYnF6yPJgyWlpvT6BPbOJ9j0mAiR/w6uzyyj75hoXISZaKF46S
tGYdTKUhWFw+1/D9y/zzbz/RIz/oAGgwP4oZnUdWARJUxm/PjTgEpkq4s5QK/QPp
X6G1oDUIhDKQ4Ug6u/kXXF8vfzmhF8g24mAdakRMpjP3/QjZKJaA092fipO1z/3J
GG7VCYRQYpDnC1Dm7dMO2Yqn0RZACFGJA61zgxYZdxoeUpYwi3y1WX1W+tnKGcNC
/sFxJNPUh8rVu0qHv+2CWm0Olv4F9XpJQ/rmUS489jxJkm9u5oD2CY+t7obw1JtF
p0MKHOccis9AjYx+ipTFUY5sgiWKK9vq2zkyyJii+mrjRYrAH13vOyvcbmZOXfe5
90aO00MqaeAbwaf8v8iH8RPsedVOvSvuaXq/+hBwDEVjugo8a8pg3KdmPSBvMK6D
uU5Q+ttdSFVrRH2yu2xaZM3mSVb71sBLOOvF8YsOo8FipUDxQYx0AeiotSZRQdVb
3vKfwk5iJZ+MqhU8l0EGykd5jKTz9VEerHf1F08IIM0LSpj0gLi9d2dkjn+43ymD
KanUxiqe30YzHLCdnviG/Muv1w6xgwaCDyAUsGxJ2y4OiZ4WcDT3Cc/0AZw+KL+7
3SCzp5emSR7k0U3VsOrNYrPRQ2/aUXn2Yu4GCCGAPElR/KUZu+Awm0HYFEImW2p4
ZKhrh4BGdWr7C3Yu1F80k1UmDFuJPXTxiMoRdpS/V5DZPK68Pnm4stiqHTAaHP0L
wYyjLjrCZ8QLedB9UGZ8XE7jpayntqUKz+sEGf3m+cfa0p2KTALpKhzguNHTedA4
L1fL0nzY8OO6qU1MXvOg2VNztY/lKE8I2zEIswrGEFqrLakQPyQFMqbf/yiUwzq2
jnRKy+JR5zvMdzPXjGHqnCTU8anmlkhBtA8VoAibDJ4olV04J/w3nmov0BhPbBSY
7JvPCt+zNQ3TeeQcwygGpgrIXoAAzcza19mHMKFwZFYlwstVab9fVUP+fSE1AVeW
S3A+MSPy2EucbFK4BaoaWxLfg982rAoVWbc9UucQ+7k4KkPSLC2jApAEArXVh2XS
iE8ZEvQ9/fvILe6BVDPKwO3z3foIvTxvLJM8rupmbyNFs12+o/6HLDM7D4AAZFtR
uOjC3MC/vhICI6KOOCgZZJRvyodXp/C/fcp7BKe+1wsfrG6Zpe2TFhC9GvXLgFU9
UAYgQK/Gh2yjFxPcIAXDqEuh6AiFCgevxzICL43LQauXIat+wrH67qCtoULMjkLF
XY3W37Fls1zvsXVLPXlDe2WED7uv264QItBuxydvqvhLIqds8hCdAyTykK1XhBz7
Eeu3Ut67piNyqwzuXoZJpxGCaek/gkDwz/zc+65VP3jMOoscvxyRVfGXQA+SYO7J
nLiOwZtBEnkjDSSzHvf2Ww6KsLvB0sHACOrbZ9rrZXNNYL6Sw9cUyCESpI7+nQ97
W6XxsUIismlWzfvYLLi57ESjj9jWf+fkU3nMn7QEpgIelMGmdIBtfPPHPKcdcme0
udwp3cxVVEbecJq/zHENsEK54sPX+LzJUXXQ0XS3+tK+nco2pSxhyp5dp6Vkvwmp
HDHyU7gbM/HSBywSA7eSvi8vrxhQVnl0F1hlcqMLrfrIlMk1HkA17CJIsg/XXdol
Et4LObgSQUOWHItUeGs4C75T8reNAXeAOrWhQZD8/NSwAV1eaTq4mQ4d8GpwsKOM
LGZSq7y5xSApPISL+cSHyHvneqbYVwkbC3bf/S7FS1IZoPS187epFrhnmTVBrIV/
3L2msrZVRkpRztpGF4cJJiuhWH/8tVjtlEbcqq9i0sGiL2u/CipJQ0q799opHLuh
85dJHpvGEumn1vYYGGtUrV+lj2EmiqLiVZGFqTwMYgyvL4AXkUPy9x54yHsH+Sgg
vSmKbBMmaR1diAnNfvWVr+C/YtpAiBSig4qfMPNY1KiGMD4StsyxosVqEbieY6+B
T634WgJzFZ4s/Bu1OUhOAZmc3izuVQ+4jEO9/UK5Lt1seuxVIrif5jZbIYk87vdF
SY+EqyOcf+xvtWok1D3I++wXXleuJhDKBqfLsFz9OyzYq10EfqD9QOK957PogwXp
q72OW2SoyO0VcdiruIQRm6yN4BYlR6rYFWp8ebyXSV8n8JhVcsGwf85msuGabDNi
a63GsmZmFX/WadS18HGosgih6sVUV4JdAoQdi+HuF0M7QbrRDvRIYiICBsr64mgJ
9IR53ICcCWVxigtJT0yZ1+JQr1k5Xce8vG7Sgf/QeX6qMkqb2ZygmdaWxQRno68Q
wo1MXRECdbphHRjp1nntbJSH9+Wj3tlrC7zxrWPY9gUGGJWYBj6tboGIWjCxWJQJ
a8te3OUI4zOgxa4rhaod4ZOh6Ff5e5HsM8JIG3w5RP2cnzhaNeCMIAzW5qeZWw58
41D3GYpCCvLmeAyMg4Dnqfy7VOURVhNCwCyV9VNBR0AhcoPhI2FfnyKHdLE6Fg4V
E4//CG9h6kjzMu5TqxFGtbta0Y1WhSXMcdqgaXmzLTNSu9tUTvWvYLte7bk/aaDy
q8xVVOvYtMUVEWw92l9SplafV2ySzPsoEg451g+YQRFdY6YSvYHgTqvIW8IBK64v
WyJWvTVWKJiO3wkbL2Cl3z2iT/jhe0BUQPsxmgPRl8B6l6WvPIujCgDdOvq80Utl
pXotYullx1vuzMsevyc7T5zYSV1rVLTjmVXmLJuDOp0Jw3UkXcN0LdACXuHthYK7
Ru70k9qYWdz4JFrZvP/xM/CV0ob0/TBR/FHZOI0Wt25MQSPjpqsd+yeTgHJoVMO6
bWfHNaOU+e32McytvaWl4q0F6QCMW5HhRF3bz8Amx7L5CUx/q6pm8TJup0fvlznC
lgrRkTRe+Q9rsQAMbmQVR6ANI3s/+I0fWBHyOIHhtEtJYCWLlpvEY2xY3qPoDGsK
Wa0VASLuDCAOE+pQypRLcE3VLMfpSyd9piJWUniBM0wTDOdaumZq5srWl3onVcts
OaxNJ1268WNrLY1tily638HZ1RRpSAuiSW4RWrBfuO4+Epa0aOqYh1+lYsHeYFrO
f/zDrbT8GQPip8/k8R79mwYHQd6EmjD4hytOSed8BySfNlM051qGdS5thU9uxPqG
HmvSE22H6kA2rSLXtUZwkoKs7q1aHIw9qFNVcs1NLoA64+im+DQyGXVyJ8h7/SpW
Vp5TZWY5/h93LluNQj9PPiA1lnZbLm4OHXpAUvl3TlMQJCuL7Gm1A9aXIMKvUStM
0Ya0YvW4EDBxArQBdsqDCBcQZZ0qNI6W+c32AxDB2mAOM2ePzzMg+cG1/TYYSF3g
tWmqhlQkmXcrTv2jUmucyP2VmuCHTO9RgdwyutJ6hp2s2w6k99ixL9IdTLuUkF6U
fjGDT4Ihr3zEupb7lAJUFUPjRTAPKHo+XXVc4BkXzWHTHp81HJztF4REUBdtl8HP
QUvfvdpICsluTR7mOyqkMmMB/VphU9rNQry2mI89ioAhaKZRtAxg+IMCg23X+NzD
U6TPGk6z3VpQzpn4njTqlWEz2z9vDvpRBI8btOSfQ57aRJwML+9Ex9JNClWBmuhE
RsJz0QrsakwR9P0pFpxJbaO9LxVyX7ifjv7iR8kJePJ4ofRnUT03WWXM/fwt93Wl
wZkEq8pkUFz1pdoVo6qpPFJ/HXSM7BQ/K2Ixnd+6ykTlRCMCU3zSOIcD/6lJQqO2
dn5ayMSpBlxeAcAafsNH65SDX8EGjWw8OOvkg6mdMKFG+4eZtIerd+S8yb3w9RSb
FHE36Y0rXF7COlG8BJ/IWcSGs9bBBzH62LWtKEaASIJym0J0Z8z9v0fN6Sp6TmmP
ee9w55hsKO7AZSxBWz48UDMl9Uc0oz+aR8r1a/YOjUaAQVE2r8WdJI7CTOB/xe+I
hdM5Cw5DR4rD6dgQ27U3D65JBhHv8EKcA8GXzo6/lkrq3FZZ81DCUmEWP8yw0Vcz
VCPxpWyG/dM+J1R7HegKizx6HEjpnXUC6Jn8HVS6XN3W6qO5WijCwSvcL1QaAU+u
pufTKCuykZrOYwcjOr9DZLIEzcOe8xDZf31miw0+xvvK7meUMhFOYHA8QUNyXY56
bzPDqGKU4+LANjZo9j2+mTu7GRzPwkNW9tkMGsVIQlAH48vTiXuRgFG6FOkguqfW
0DxauOanIdRErqU4rTF4eD3rmxnlmzZ/iEdcU9+Klt41bWBd+SaugoRfchu/qBaJ
ZIw8uyZHkaUUzvMJzAiOGHvoVAliCy8bsi9q+B/t5RtUHkWK2GNJwE7Ps2L/DZ+e
oLyt1kaO9c4l8wlpSFcbBKg78wVNnzfcBxzDS5qxTyMxrje4c9LsRQktsuJQHOCW
E2lSTsU2SIPqSKvtdH2qkVTwl2vX/z1U/K5u3CRm+7ZCRHFvK1Jy+mIcSpBv5msL
CR3Lg/LBAt2IAULIdrlA6zQLox0+O1j1EBrxKDfKAjOSjd51Ray2MjatUVqS8iIS
jLMZaLyBBMZOt6POFc2HpExO+KDMN9Ad9Ryfw6nclS8oLytATLPXdHDDFRvHmRql
QtJzFOQlGwbxLPwMvAaWqwQvBbvIo/6o812zJISnHyb2zE536e7NNFFfJ72sFWpa
yEJB/UvneIVaSkF509DTbwukHvindURyLAxcV8dMbT5zjlUlLftsb4jxhOjgfkG8
it6mLzBqWRvsWIzUALP55VizU4JMoix6mE2RXEkPFGQtTEP1HKwK0TZggOKHD6Ck
fEogqQXFrZN/23iXT7y/13Snp/+UPIXaMWnAK5L7NhxAx3O3/u3mrhQBsR7B89mY
p9ZAswr+gqCAsALYCKpblLOxOBgYTQ6gMxCOtMVh6tZNXYI3CbOasFAujDE+gQ8A
PXTc25f1S/Ej1U1ELlrZ/FAqxT/ZVWNKQPOWF+X6wuRVLMCWphhRVXoPWg/O6A85
lDpGHOoE7UnkwtSx8/bqmm3Iuy3LQm/ORHMlaZqixg5yMTkAGjw0R5i+FRKg8qYH
z4pZS9rbQzAwyqjIy6cWyJvMNeymfC/3fAb0I6nf8r53XkkAs5jW9meJ269HNxJ0
PNBSksLqxpW3S5WET9MRPeKTpCi991Kwb77NSPiZyLkQT60V/MafPvO3IEyM/QjJ
IdK9vDLMrkwCLxzUH0jR94ZpIdMeJCTP5xDm0vqMh7tNJkJP5Z2K+r1m3c8SaWEm
uqpw4w6W3FFU0q2Vz7nqFT9suo9Zr098332RPJvRAP07pyWft9CWncYQ4NMeuFAY
OUAXBhikN/vbuj+1H6gwXP9bwRB8i5tKKMG6BWdYEdwNBQ3cg7OFJySe7+lGtqhe
Ki/ZnGrvIZ8Egfa3owwccV7Werw4eDBbAzoTNZK89t8y00yqoBcn/QdLJUeyl/ea
WGPLw4mYMyd8KqpITOsYKRMVBXey+mYl5Bj/17d3ZJrui7drTUA18ZIZO/2IAKMs
yLl7wSBkCZyWKmlSCenx8goMIlrJPYh0ldJT0qfcGDz72oU10lv56igrs6+f9dt9
6Kcls4LkA5p9d9zVbKM5MfLl4c0ierKdaFzm8fnGMvuM+2KzwBv5S2wK2Kt296eC
119PCbYx1W3scksh1KZl5TPnX8H860jDKw6PsnyEBQBZk6Pj2tDIxnNkT9JZj20Q
J7dnfLSyX+kAEhNHAawD9GU9bGufySzoo6QkFULUFsFXYPOzHOgc26+Z+UHhRwEb
nmWls5uOUB2ii+OA3KEss6gy2bpoQ+1rBm1ixb6tLgc2ayKR3ika8v4f8459S2JK
jals/noPI36ki/t1DRCWgBbFKyK6gKmIimHZYrLYbkBS4hwToECxS6bo7rfqmm5S
q3PvzantzT9Wi858uOfnQhoN8uN9faBAsndVQQvw9SqaQ+SVrPpKxh4f4Gf0SkdC
MW+zk/Mczu4RP50zgf99YXyURmoh04dwl6slwQ2g1P2thr05YwESrvy/Ks+Mh/ui
bXf1KJhLg893a5t/HyEEPC+6hHaAfRfCvMhl9ks685WrbagJhnsoarj324stR9Wx
Q9ukUlglsqp0EsXb2jaH1DCQ6nAfYgwoWTrXTYeraGh18edKafiSWCVI/d05aThZ
mdRajYNHfmysti+126+zz/0ygufksfo5T1rdUDJ205Ekxc/PNpBME015Jy8pT0Xr
Nd69BKr0fb+c3bcJJrpoOkaMUA4r9J7Hq/FSFbOfYNMcrD0Ek7sU1rASMojZruHg
GKNt0m0BELzU3InTEBWrGqVkcYQtxSopM8vGxsa2549K3RnLKcoHlOjvPhOuEz9y
LdypAq5H5jL5pq0mZAvO3aMlbHDDNvY5dTY5XwMP1KmDHsqWvu3s58yrMrBDHg1x
Gtz+5wIY3wndfQlWR7krws8FM67AQsfAmFd/CuPaYAqqSYCIb8mqaE0bU6mB3dHR
kylgQx12LE9CIL9AYA2b0GaNmLSWbUx9pJEvFxsWdIdIAsVmMhqeZAHQMlmwuARC
5PnCxHBsWXmUZVwnEY0d0ym5pG1yGqZ4nwzHm1m89gPUE+IAAYJ79Wsu1iiWLKf3
hk6OIgSHIKApOmTckS0DXUlkJPzzqCRTCqx4Z6laN/n+Sip8hpQ6bOrljg70/JpN
tLkqThT7aH91CVT2LNp9Qawq1NwflaYnTuGPf3Afm7+HwtWfeLWUf3k77c8zZtvI
anlrNHA7ZaTRsVF9YNnvbcZIGkxsShL0YxZxm6kPMRprIixfG1LOBllfBXGx30u+
bUuPH9+rrRUuRhZm8jtlUBvG1E2V7iSv/Mvw9iFlpIE+kK/YmzF/GgCU2WfC8OVa
o8K1i8h6/H1XDVp7XQn4QPnY6NRxiWZcm0Nrobmq3K3N2OFZ2K7b/nt33ZvBYDVB
mvzlkZG07d1d88QzF/q5XiSI/qwZO+yPhwIoSW602NapDjVh2sUvgHgzkWxgfouH
QvClVCGraj5Hs7ISt9D/DvP+nzJFXFIIX2Jm28RuOo39Cn+Jiv7MMD+c5m2/TEzh
UtkAsM5ybPyKX6ND8NN79ffr2eXMRSlqTzhlMA8wueMOg7Ra9k5jf0eqZB010uwd
NyG6SOMJLtpDPtha+KqDj5wmaii51UZfFP/KonzpAND1d5a5m9XwQHUbBqXG/qoY
aconDOauky/VQy9GM72MBGD9FvRxL2HtrBtoweYb+BDmczprNlBmm6CERpXDj3Ly
zxvkTsdpFzHypCjPmBt66pXOrzdbhjmG4lseVptUILIA0Zc7o6v2/dOIJ22KNgW6
Y2vdC99KYyU023Hq4IJS/uBNqYWDO1vuTWz2QvJGrJ6cU3jhxROL8zXT1a63u0jz
OTRD5/NSnh5iQFYTcsixDAHvC6Kk/oe85CeeBYGxkVXhG4oJrJYpCUPXP9JeavYs
DUyI8bUZfZepW5APB2wRqxCnPSNWATzfWvEC/NIH7yO8ztNT16hUN0vPuwwv7JrE
SiY8tBOukKYSwysd8PU3p508A67Za+j4r7sOu9LMkkkFEnnFi3K9QER1Dqm0A75z
RP8DTWio9S3KPHgeobXGGfBs+7CNrJc2y5cPuz/qwsgdwWKxPIlAEieWcQ6aZ4uf
QTuaKzwxcbe1Tp5z2X13xt9CBmiP8QNFCIScn+JxqopWSEeWcyd+gTpglFjCyDUS
O6mOLRT29TK9krhdz4B6jsWFVwy5h0u6CFWg70mn432PGsyPTbO4Cl8IrQ3DkTOV
GeuffjleiBzE8XcgQ/qCPBXxWQoxbpZVhs4JI929JWQ6fCQYhAneeU+I+ludwRRz
udZItIZ+igLdx8nUSimF8ZDQYui4vUh/V9PElWUTxyPynPw0XvJ/2OZ4NKicHQ9m
/RFOJLV8RbCnYhgJycVPdBIVncbrg3XZ65syQNhA4PZgAbXbiGeMIehmcQbJHUJG
0AWbU8wVXclnZoH9DPzWUqWHBMk8xC1LeR9/xTuKOOaA2lMbrNhIqPmRt7uactWG
9P6KxSPuAmsGFgukq3A3zxdka2WQ1WFm7kUPZie+Grvw6C4gik0dkIGNW0SOFfk1
sUUgCCc+kZfvxsjnh3fmw6EXthUYU1wQLVfZRimNXzMzNsjPH8hIvYH00l3AAqcy
vozkxv0qU67JKlCrtAVQqa4Vk/btSlRHXyS2F/za/vSa3raEB+nOHxkHrB1ypppc
wSRkk4qiHu9zH6Xjyz75tT1DN0Tk7DyC+bx+VCFxF6wALs2RTz3u2qY4JCliNHhd
FUR2BpiUlBaagdGsxQwif0ELfjrpfoMCjN6obrTwgwesSiR3ijp3uD+FpnWnT9Hz
pp5rFsIefIAD/1vhcvVovaovAyqeDRWgY5tJGF3CA86oqeMRlOjT0WuJLaHrBPM3
p61NNRueUBIpx5rd+sx9p0Z0rY+Ios6CD5hDNXpFx127NtgWwqT5wJKb4ZvF/J0G
TDtHvPcHB3WDxnwHy7WBcGLzMLkhv+VFpFaqmMnH5U6wWIYlNNEJMj3a9u3mdItw
BLvF0a1LrC+ysQ67YRmggVn8SXIHJ055W118AsLnOS5wmNx3AEfRWKBDxN1AWAnG
cxKgrxag9z6B/pktCR1zEyLlD3o1pmwMylmuIIOD2j0uk/RbhKQukLlPBcxD4ADR
gVfc9nb8QDZqg1Gn/UDiaD3yDdxBAT0gFyLFHXStqk6YTF1K92zWFF7WZmK6zGuR
1OOQOz9O8Mp/ZjntTbAmjH7mdoaSQkgm1mUCiTR50dz8hiljDYWIIT0UUk2FUMab
NoAvPqO5r3VVIBPmJae/l3NlDmdaNXIMbSqCLsOEKlikYt6awo/Vk8Smhr4tsfxY
AP+mM5YXeE74+6ZrYD4gsQWkaXlG61BdzlIIooYMjN75bteeLZ1aeq5nWylJgrlR
8inhvuDj7jL0nP40wZxX2Hyx82v4LNq2YecAun9JQQFgWUbz/VD0EnYAvpD4WPUT
lNdSni1DuhH/z9VgQmP9fBUK595RLy/ArxX6sEZczozWR8+bpasghT7Y2pQAbmlz
XMXRnNvZpV8DNQhZxMpha+VFQsgR/IMPmJMOHIkdS8r91vw8o17Feq0WF9mRYuun
0lX0+rqT+no+79zoSdaupA2+xNqTwy6Xt0PA24YAZZTQK/663FaZb9SSy+cQ+oTg
vxakxYSKB2vlY/XXe39EzA+QATU8ebNCIPTu6GwHGw6NR4LjYqvUFMRwkRiws3tw
SQehI2XCgCqK3R4wMp4gQ4SJGHawcqG0kSLM8FTt9Bi/dOdhTyjFYD+I/m0XygP5
1xdbtxNz/t12CTQOmffOAfwJBiFi9sG7+hr2N+eL0r9Z/ZrPFtCApJUqx9U8+lZZ
gslb9C06Xh4hz+h9OmkQ+xxtq2I4vYvyQ0k95yG4DCsLBlwuRb90jWz0/5AIh20I
prNxVjacf4PUginaSY2D8Y+33fw0qqjWtibBOI2zFFyQJetgKpZjE5p9pPmBDj9Y
bx+/9+cIZId5Kt0K4BJSVvy5+HoGKKnl3R2J1/9MKexGTJRxby7qbAFvfdOl3BiL
7UdGbwzy3Vnwh1+3faCEVg0ghhH4eYdjHkYmnq+dIbyXwms8uar7QDPHNRYnUvDt
cUUDtM0mVGt06JXxkK3rn0BEYl/pBUw4acOAsSTOrADMs2cphcYAeleI72Zhwwp3
BvQFinkXy0+Qt8v1iFsLyzEFiMRtGvy4k53AMVww6g0w5+51lZje7Tu6oqh/QvWQ
9IRlzIAMRF2AGqX1Z8Z5JyhGD2k4hVZiqDjKkWcuGhUd6iO04QAo3gSIxUbHOWni
iOVIaXE1GFajVsB51C0mVWmfuki6lxsbtO9+X7UGcb0O31JJgD4m7Neyy6mmvDMj
jTbcTNBOMHu/v2H0YPidEyMoLETqdtcTH+iYMOdhn7U6hVvYkLOBYRSvRTodVwDt
egsdV1JJUKG7qvMX+XY9NA8s3HQIgjBQnqk7Qhs9UwgUwZ2k7XomiFS65JLGykKd
DyUsFviCMABugIA3mI32lstke5B1Omm3QMEZ0bD8dIcgKS5P5HuZ501eL+LZb4g1
fbrruzWlEN0/BHNmono9JMBjyUQvHRYF1b2042b4LkSCy4ah/a6NOrjOpXa4WLa3
gdULC6qeZic2UUgYXCrnNpdJywiefCuKZqRIXBFitw+N1n4I0ITwCWBvURKgCSkT
3wc3geRdmA8jKDN5v+da3BqQkM9/5qSZNkU57Xk+ffPX93u51ggvWrW7ontrF0nQ
4e15JQFfPjh/BZqpUX/rd98BsEhCjsvs5A8vfX2WEBG7wZkCPw+/sQuckpDb3b3Y
+XkC8s3vrf16TFzdaWQYxAJyqiTnM75rWiRi+GpgIcsfTcT2d9WR7Mo55fngMdhe
lvt165DajVmuYyGq5pFKkpQ74b5/tad0iOTi+fqDqu5BXqoH6jYQUElSz+5QM1hc
uBszZA1M8MGaqAJAm4Bnxv0lZ/xjvEvn7Alt6kjf7CDfFz5J8eQnvr0S7ZASHTBE
J3uwxtciU5Xrc/dVuisDcLf7dODuc1BMLfUVE8PaE3TjMwo3YrAygvHaz7ulwdzX
QJLCqxthOFE+EpaV6SNweNoZrbNBR+S7swcXSvDWIZ5kSCwa7jRv57ODzr0uqcxz
OGu2DYiCzXLQr7V0ilG5ryoDFkuG0pe+e51qUwlT8IhbGBbuynG5oWfi67kkgXwE
eAvKYY+dsK3EeGvRVkGc9QkHcOa0y7gA3cXHh+Ura1H10mKAkiA2OBP8RRiTUZcG
zyEpt8gJqpreOQRgZSxt5eKlJ8Og8y0hEHpoLpclYKdp6SvNGV1mX5u8vVOHmzXZ
tcKo3M5oaVo3DU5hSjKviAjXT/MQZWrRO3xj97XuEzNDKwMbKcE0Q6GXaBAVXNOS
EYtPuL5I/hhg5EzG07bdWGRf8ZmGDb6QQXGzcH7k59nfT2HqG32DwGUjdL/nf6Xd
ooiw01IuTV4f8YkAvP5ZpucTBsuy1YZBKg9HLIU3lTtV7rsvZzaUdTd9W+6sesxo
j++KUJf0dpwrSvMlxPC4VSOtbrNvxCM1OPUe1MjXngnkcE3jJ77ttp9sr5Kqe28Z
W8pEKB48HHPr/kd2xCXks7GqPicyOjR1tAhvN+WhbMCYBajeqTlQEdn196I4HIUN
XcC+NuqEBYzn4ynihLzMBiJt2xy2XBskJteCnzkgpMmB+y8GSO1442KU222We+x1
kQm9Q2CsUYfBS2hFGUztMcFGfUT1lCH8CbOZsO2GlJJBlcrNSgz41VAuAXmmJ+Dy
GvdsTL844ZLDbIthV9QghPcwlLfY0JmNEM5JMOwU+mVDNocD1eHKaJIo6DD7HZjR
IItk5XKN9faGzo0Q3L0n5ZmdvW6+uvbJvUFAdBpOpm9ETGeryhtiFuuoCjsSIjcl
Sb3WbJUxG0dYZ/Yu/y4eMvbiIDZk4QZDKZyGchjcC03uuRxQ7iZTeHSdpWEre+BB
QjCLj6696rJW8dhDrG25bd2wnHIdrDEcPp9j50Ux22dOso5th2rHWsa2KH0OUfR+
MbuN39FMO5CxE24jYSkCxFaODw8hMoPoMRdjVEds8pxSDxhEw6mAgJDNTkdmcRqG
XEt7c67sb0tMpdogEteKxHbrezywpln7dyvCXkvS0Bo/ZFrrdwy7HvWxMHr17Uh2
z5l/XFiyGhkKtyrV0t6VXt6ht6fuc4rKtLNMVm0rCtgJVWUd5A0sjoToqGUz7f6W
/Ep7n/5p9Y5sZuCz+UztOmYGkxLHOOY9ujoB+DIx3+pKsc4qZ0Ia2Opd3DPiQnC1
+ivuKMQrc/7yS1+o6rf8VWNfNKwKaiqVQalK0WFEi3Mw3NnfJLiMbkHlcJBkAXSb
I5CMINpXmauXpHZeMYrfMWOnt1kn6JLT2a/v7GEnGMyPv79QoKBwSZpQ62prmbpB
4R6J6gBHxmgZ6hPh7FO5nqcj+d8pMb/sFjOzBQb41QSoZxtOhKRitQq1qRMpinc3
gfHa463BZzfSOT12jBQ49Vx2gUtYRplAG8ARnPqWwncZWcIFTPpZe5USBQpkwRMB
URjBNKgS3LwKcqpu/IcYZjVz1ED4IGjl7P3oa9lujNeeDktV78S8bJJSZVRpmv1s
qcRo6b97rCO9yTTxLMsOKTeECaaw+iJhh5A8MVwVrhFtKqQa0r32FAiYYUZoscEH
6hwVmZGJV7o1Iw38FJbA8DvdbsJYhGnFDFcVVtGgNGGPiyOSPMMFB2fmTk9knNkx
sOqo8fjZE0z0+JRrjnt8wjNpfWFFwbBUO+USVY9TfBOlSak6QOzpYJTkDHGzhzfl
1rR30FY/fS/F+y5r5OvR+dUnpoC9IDWWB+VyhQQPwHhdySSt/Hz3D8Tgnk6ZjJSR
p9lP0pzVbkzGcTPX/mRk6PDYiaITHjTZzpYBW66AKNdfHAmXpuoW/CX4QwkzKcL1
HgrJEbuSJn9uDuDs5UIdnKlaQkFviuLOqP/8ZOACJZnRKobrCkrqbPR43iQVF+iB
IO509apTzxW7MZ5Q8lL4z/WcokhKMRhOy6x7N+PCtB24UxNB92WUHj5mIQFpenIv
PsgdDN7C8XxC5VKhQ+hbPBuZvMXhHQSlb/Hnrn+b4ZJ+mkzk9jTh0depkXvgpL1I
V+0lKWjcVMTOpYZ4jorMEYuttYQHFsVqKB5Tm8i+OPByHU/q8AejEVzqzQYAbTep
m1SkQMbE6WCWuxixvQxU3Oa0T/OuQdtHRLDC7dDg5w/ZpH/2PoU1aoFU8UW+Vxkb
8TWPnaRtmK6KhGu75RadocNtlCxkkxICXgG0T+iYo8cIo+iaUThXXtaYxdsWjfF8
/B7taVvYGIMifPo53dwmqIGVSGNVseSV8IfBKq43TZA9fvpxk8Y5OAmZxu5dzAyU
XlgQ/bVvEB2Gi6/+88wNcaNVeJhgA34almLm1aHwDPZBDBB8f6DqwU61/mFAiI92
sClCNPstB0xGqdxrKM9cyKkmZJxOX8jKecPl/ur0AQ/ububKVAeuKqeeimTVK9iS
s10NoD/G8BaW2ebtRp+L8g5zoB97ASc9dAIsPPlNzg9qMq0hwD19XxymkYUDxhK2
dLRoYclrsGZZErXDuUkxlmWr1JFnxuTuK2PchBfq/dY9WDeQ3jHVVEfySqplzMbL
yz4Ho99Z7UwFPCuu2mjUwPW9sxOL2Ei4YvyYaJLGwFIRPEoT6EoXofbKmvaIFuAj
I61tR1mNYYfYr01lgn7ekRuPZy/P+d3FtnS6NBLqcfr4j8H2jescbabgQx1++Cx6
UygrNP9Z2yVeLwVED+KpJna0ouX6uaWggz7XMCrc/CcRxrO0pothis/BlBGWpSZU
pUF5d3oRn+IrAPmDxr/syuEsBuAXH26mUyw6LczwajZO/gs5++nUFbiHTeM8N81r
+nQi5+axCVRKjlJ06oKWA0DoTn51Ut3eVqFM8gSi3KJiXA5ajkI2k/cmdpbc7n1P
IZHMqtJTf2u6BBG2mU3e6/nOfj9aYaP7UkvZx5XRF5NLB+CeNBsgW3IWsyzpeMcK
L+JLHXySHLk9NqK2p5/tIWuIjiH5OohbKDXg/EYTEsWU2KtO74DVjmPuSRFzaaqc
fR157MQygYP3eTxzxgWUce79gvNEALURx4xb9KodZpHGCPVQSy9JPOUtCmLB0f27
4HN0pCJzJRWIHf4otcn7WNe0wCnQiD7IxqAE3kJ0dTDlYgqOMwNV1Au5OuhaIw27
JaDbBIQqU8suiwo9q4ozSejPM07wJ71iifbne/IEJpFPaecfbJ+dJG30earqBwk8
UkdRF2i2a6cgVi1eH5ZJhS5QbdFM940B7ICxRz0Z3zJAONsRb6ffDzCQapbZ2RI9
kaB3Rz2e76QDlO11OAuOWw4Lbuvgpl5IlQzGuAlE8VfGW7Nmf2ua4nWOp5KeYHng
Ro/UZspWHSLcnsSqwBZuz4wDFzs5sTfqQEF+TEIGGBAAuJY1vQQ4qfvf164imCBm
lCXJ3e0NmFajwR0a3i14xNG0ahvJFJ/7j6LttM18IMLBuNDRINh+7gz04HIsb50w
5aS/7x0epg/a52oLUGszyfBAv9geQMyZEJxo6IgJdG44KsBOAOQwZYQw/zEECwos
QzzLuR0dzKmyUlzt3FDUwuf5BSal2KXKqzmnLb2e0f8/JU81IsluwSVTWmtk4u3i
rC3KMJRkJgb0iEpL2FoNwLbvfIgHcRITOzeMctjzs4VbZY6f9sI3vrH0qMxR7lFC
hFjvdGgt2wo9FrfZNuc6bjZsabwHl0w/LcEfB4gItHX5C0P9aQhkjFAPIMMd/Gz9
X0llWgDvMu/Xqt8CB7ZnR8pGEXrx+yawLuHyihwOSnDUqqVBbydapc8g+KBx3Id/
5JapqbJ5R/JnEXFxffZ9cz97IBtrcw6fottvbhEzKjFegVnRlPuegIibOl4FsUpG
M7lgzlaKhCxoH+rzLB5KW5PlVgvIv42GQTTX29FPjdKU9Wf4oaaeLf4HWxpZ9mEu
va4eagCUwcS//eMEgJmuQzFwc22ze2nyLfP2OiYOdJHj9db6pKlMST6nWAMCgzV4
EIHDdjr+JnRSJRFp0LDAlwk17K+56KEkGou2569lbDPk3G/ORB1VY/BgECUYqjvV
s/d1aESBJ1oX/kqYjo+51U73HCvssdbVdzi5Fz7uGr9H7RVHU6WrOlW13LNZrm/7
IKo7XC7vy8zwZwc4LNx8VC7kQXsu7Z1TilaJLO1CZDve3X/wvsX76vhAOaHdxl1f
Bn+KSXVjzC3hVvnqbTEbbpSUQ7EvMbj8tyTETZY9LW/NluuwM3yj8XQgyQUVwj94
A7E75THSj9+ZsJc6Ik93+op27dAdc5nIu44/9mJTllxZgua3aV2UlFUJBNm1nN8x
FeHcYoKnzRAxZJhi32YWicKIG2pLDiN29QiEqgh4kLBeCkgaUjwe7H4XBJOoPaos
MGtQa1QSQx94R5NRybFgK2n6t1q8Qd5a9Gv2i2MV4ZAZfItcB6gcRjnsJwpC16u6
Lg6FHIj68bzg1NG7XoA+UQB2IbMQWVbJEbxoc+TbkpTuGFV5a0guz5k7gP1qcbud
XX9E33zW1UJzmKx54ITkj+1vT3jVQs5TdWyvIhGXTyh1lgxxntgKfflp6HLCUV3E
L2QcwvNre7ybcSmUCiMz2uSCOx3GpM2oQRLqBJAQzZYVQ969+SHcwnh8JG/qAWfc
Xp8goTKNAa2jVl3PNum4Mk0PUYTiyBfnDqF9EPTWt5xK8RgEcvGXTQGJuv03QWYF
x7hQNifSZWE0NzWCFgr1tir3ygQ+AQp5lUdTtEGV69syjfCF0+4z+590JXU2SKWG
TzuxpAVy6RJz2We4t4x1GzZXTCPmgy1YAE2FKejrNwRh6GMEvMsf7WXjC7HOb11g
C4/+b57ebK97tAqwDsCBj0hMrsMD8eN8grAp3cv8fZ7a582GQ2IGXkeqqMzXRcbS
00VUEl/M1cbcUvB0xlTveSA9Cl/Y+quB3eXgkrpqD4rjK/8tDuEMJHmIDG00QRNE
gRl0V3lUhf2hsKJtfLOflz7BnP7f4NhgJDU05vHWPUL40w/fcUdUaP3+Z82BHNd6
MYEPXWvfvwV+5xNIiFvR07EV52pUuZLwdDdtbg3gvL5uT8ZiN4RGGF9cgAl5CpOi
8BPxLgsGe8XgNTtLqBvAlMnWQCBp3hmVYTfv/RDCjZNi+RMC7YIovEdZDzP/eDf7
SpCXD2jM8cfPRWHpjBiJVUOy0G1615tpXO3/tzF77JEth30cb370Guah6o3s+Vor
xpyiourwpgOde6PELM+qgo5AQDFH/qxOe1GJ3qTHQSYMgieVH2cleJA8ysiPPpX0
lqNBtqMeCCV7TNQj6OHNLXQ4s2BPRd4GqD84VqXdkTHBLbB6J8nIua+flzdzqD2p
KNHjQSGeVaDMRRRo0kgF0/25HC0vC9+10OE97cMfSD7XKf57YBrJMURcUEQ7lTNF
5+cxxrtWi2/sWpw5fnVSj7P3VO9EgbyVZFKBlYLlj9RFRTjr401Z9dmhX7bWjKgc
pXk32M9oOup4SlAdes3PnFfVjXrx+6r/RempHyATMCFJ1Jo6vMfwVshICE8F8p+X
ILNW53e9gvUx5j+DJf5pPlP+ofdbNmahIdU+ccoj1XXHwqUeMUSTyrsscjD+fjYa
b5vhb6S3Tv5P4Ei2nS3uFcg6hERaxJrIuL+c96LvFt5BaEaU/QRO3v2M7GKuNJCh
taM+UMg/V27uY3W6NdYMlasyKuWWAMMTK1H5tMOv1t129ijYjY72x6pltNvuSMww
K+Ven16blyKPpce/mqQefHu0c8l1VlT98FF5RX0OQQ4M5/JozuXiqMpcoTfrJOOD
DeVZ3Fv86oof3uW9BRLuTgnyqAfNyodA2b6pjWYahat6gF7vcnnCLvby6glq/xb4
hP2GCtv2knppKaUcZO8uQKi2/NixzI80Ul01BZDWjhQ4JcmSnFUwdwutD2PbNTiB
Tjbr4LtVSJxSSKMDQk5ncJ1Z/92WH8t+IWm/Opwdk4xFl3Y9kTBUCOWB74RIf2EE
j7v2T/tOEXDOPy6Ve2AgsrEwfdXutdkqxaaL5DMRReD8Bnq+Ut9qAdtW+RS6MW4l
6Pc268A4sHRi9G2OTyKiJkmyC2j3/vfGaNnwzowFumMngMX/zcKnuEI5tGvqQKst
auh5yDc2bZRi3oUItILxCbxhD92gCnCs5irwie3ZNTzBCRqNCvuDkWqawzQsKAd6
0td25t8rctZKcQok9Q8qUM0DMPcwC30e9OHSTnsyUHFYdXXdbBcSMretVTtlEbk8
US8bVs6TDJf+cHHcx/vdvSgNZ1OiZhY5ktGg24R35vpqG/ZJ+bescH2mBA1Qoued
Mc6bxH9BeNR6KAb+bouXg/SUpn6B1eat9+kaAAMF+Vl+9d3wrV7UbBqL5ZAMv3+B
zliZOzkWq146ZDwnNvno9/Fjt8YFlrC9JSYrZnxyOGZu+sYqdwaJ1p7Hj157Pe6W
7Qjr0zutYGu5G+GtvaLIZIRh/sw+4gkO2gegmP2nmZYcdBfR4x3+2RrkdsVGo0zK
owXg7fPbWEdaiPXATeAM6u70HOV/slB2tPRwkpJt4+SxN2EbxU3OocgwKIXYqM/2
v5jtNV/VBkj7++JYfOyfbN+y7rSEmhdlKq4L2qtmbNioVLT2iRSEF7svJJLFsOqY
C20wd/vMGaQC3KZYwiAAib7FwoX635TfidKaL3F+313w4+FKPWBkOYWwl055w3oN
H2sToA1ZSPssepRGFtZGYgx+GbtWZ3RcyTtQe4rhYzQMvUFy3vDx2vKVnb1lr8Fc
Y5nTACMxw9bImWiAuqDqbep7H50IG1bot1GG/QHhPjkhqEG294ZVbg366zEdh9af
qqwwzBBbqDWaqH0kDn0oXAABfUJbsMv+ZVMNgTh6Cz8bDdz/IzcP+Boyf90eeGeI
k8WsxOC6oKGdabSaJu8kDH96NDraCFunyvJei+3D1HjWNuoSVN3A/s33g6oW+GE+
IvvCw6CeE+VOxlPUjMWrVlLS1c8ZotGM8m8SWcWZaC9Xkjq5CyD6/BLDAcJxHOlH
Sp+/AZmY1D0LIssBC+kTKN7rn5Bek8M4FiLl+/qLhnxH6g/82NvuHRILN+nfBNPv
dlLjg36QfJKCh70TqkMl1SqlrS8DpaIo8Qya5LbBB3e6g3QYkqpykpAKj1MKq/P+
g+vUieTmvXIdEr5HRHwzdPv/6/uBnruv1Dlpheljw40bWyiNAiueOIxlXDGBMPuT
Kp/8N4FsirEAzTRlQNwGUTZpALodk6UrlteDSToUG60HmMXuGJGjLVPM3RfZqTH4
1O9kwqjya5SJZtOyz6KAhhizS0Y9r4um1LBY+lGWnUG3eDSq3UAZU3MRpRRNhg7Z
c9cLpesErXzbwc6WXjs9a6R0F2QV1XmloSQBdh6HB97DdzsWg57dOjRMKwS/9J0U
Aygu6/1MibeVLeVL9X2nLyFnuPHjmmzO9yqyx0qD/ML6h102REGWPm1I5F2XZ5lY
nhIiiMT+sEMkRr6HfanQyDOqsnfQbFPm8yVTVKZP25oWDQGIIRbNv+qp2kGL1YnM
jshe0irCri6BWcijHgKV8cC3NSWDKo4Z5x948KQ+vO7YzZblY/apAa8zD1OSDQKz
kx+PufX/FS66xHy0cGlHTRyZGFu+pi+XJX/Z2JXRHcQiAyEcDDRIkS/qjIBdbuhF
KWWO/kFdVusu6S+c9nSeGI0YbneKwg434CAXKh9f4w64zbIItpkt8NtyGZhL53ZQ
Nhlj6F805GoHb19i0tXCBp7tBnXYTk6gXWfo1XWmTqWkEJ+7lERFEI8FHb4YhWuw
kge9ynNp+2uxumYvkTVRME6RQneaNhW5ltsVsfpBGV6tNJLvO9+EOfyOxvncPVt/
4201vciGyHZ4gvbBl1Fqi4iHPCQ0Irjhoha0hWBvy0ZbFkLulz18cBIK7hSfZIlT
hKtfXXuylhEL6/aMZtAYWFGIc9JFuCgakgIDE+RmkPYHeLC5mkjNnwrt8pYwngkO
GBc2bP+T1PBXm2HHQLk1wAblYPnOqgEaEuCPnxA2xscR+pLR+DxuLv1WvyRpiwD7
SbXef5TGUXB1PKqr3Y+949ImJCMTSHo4qDKWaoh1dQ9HWrO7DxY25Q4XZWZZV89J
bhjYAU79mT6zkH5DDrmUM2XPWe7UAlgPF3J7yU2+bpXdxJ4JMl2gtInSHMVsG2k5
ujAleW9tlZ5dRfJae3rF1dMtJfNf0KmRpeJwDaAS+loxSeDzUrGvT4tyIKHXIagU
SHPAsB6g0Dgg3SOmSkWcymUsjWHiWAiaI4XP/kw5On+NvzCr12mPfuGinZmSpxIe
xmkop3iNmSPc49DqAonjbY4V8wB9shF7l8V4gabjr8UNMHv5s6Z37pSadY7Wg/ik
8mFkhqwxr40vitl17lavDDQdBhZy34HheiW2d+U22FKaXxL952e42WIGxOAO2Pwa
q8hwZCiOQxCD5yl449dNkM9vFSjCG5nPPsKA8HLNcc68i4fXNeSRf7O9HtgUKEGE
8fxNJqp9ZYl8fUHUgiHEujQlFnm0j4VbZQohdJoJ4mzPqNbA4SqJQC8vJxZxzE9o
jdhl85hWdyKe4Nt248VJnRZyetyxn3Xw7r34Ll8p2aDVfBUlwskVuaf2r1b5GDa3
MW+SecLyWvAnYF9Diuxaeofdr72x1H3ZlA8FOmSh8YMNrHXJo7krmC6fQDdA/5Wc
iGr/fVlNVamZS5lDLcl4w9UBXTJTQeiSb0enYadYnmUqbskRM/HIKc/EYDAxvJWI
xM/Djkmih28Gl7O7h0ZvQlIFXfE9cRcA/qWQNlWIa5ncdLM+5IvDrOsW/sBLWdxI
V5AuyFFiVcmmzt385Mp1LTmxj3HPXZnpQNo2YXVCrno/A5IBfkJBKDmBBW7BXrfU
mhO4x1VINMvp72foxh+MhHXOjBG+TQZoDm9SDP5a5U0XYlrXD8GG77F596N61sE+
e2ALq5UHPSF5jzOOnU8H4LuAK8iz1jy0d4JFD//Anvxa6PL+RqWfCt5pdiWox/sL
EdZn5MFHEJOPVuU6gwD9sv1ZGD1lHMXARmku5WaJNU3fSnRJcLTz1m9yu69TFppX
0hU+S6IOX/aixZGH9FmlFeidRJA00vTvz975k6HQZFNLinq3uZm0HYWcJiLUsfXe
k6Xq89At4Q5FWwt8756IefgFE1eqhgga8XC8Wkv56FoV9UrFivymVR4vYCYqSlnn
2aVFCSBGlRvPcAnkNUO7pafz4ri5nohSd2uBLrCFctn52oyRXqDsVy7IuC7i8d6O
q2fv7FmalgWVz5u32PiAxRFgiLlSJ+DiyW01Tty/seBIGnjJp5n6rxSRQpXBOdN1
Dn7F8MrpJFZqcyZFRBVBW/RhuPT51mF9PLkD27p/Im5qHZ6ICxGpnvKIUoJMu6yx
AeFNd042B2VqUJ9IoLrz5EcuSJz4ZCNbDNz5y1A1WJZ4r7IgP3z0RJ+pGd+fZ9Dx
Ogh2kn6SFjw42l6nKSUCCzIWMWK1AVwf1EQ2snUTaQiMIsNq4qczq5bUBAEiGy/B
n/n1Hromh+rAuMkkkx4H3ochUdSaIbjPVsI6l/+MpS6eWAv4J4ZFioDEOzg89Lic
5agy5CJ5OxUfVCdXrF2uBs2mwU5L9bGLwtsbiq5aGiegY9PYaoZ6lBgb0KRJJeFG
1w1uHbPg2BsfM3oT+MFrl+u1g+sEbzPO0xpSnvmEue8Sc85vWloNYaAZBn8407dC
n4jLmkJwdrhznJ6UPqZq8SpOHYynP8LRWbTDNWfwIXXmgky6DCQfKSuSp6tvy83b
O1MlVcPYbR0YLsgQ4iGiBXlesrWpH2J5L3HKT9hjzl6dKwTNXa8dx94DzoRslPOm
KzeHvOIJotVaLhniJ1GNDsjKXr7F5T5aPle+8P1DXA+MprkpG9sAYbOmuwNwC1Ou
OOEBVv7cApgXixniftyVULytXB5TuCMTX3sJWHkw4bQ0RiwZjuMjkLYd4KfQW4BT
ZxMpLFoqpd/IXuBn21AGPWZ+En694T2P50E9urgpgiSePTiKZMkEXvHCCfuSUBS4
ppy28AQrIMB01DrGqeqcaKILXIwI+PSU2VnXLttsiKSJ5xUpexvmJd6pz4sOUYgb
GZhnrygE1FD3bftY/QSeGAJZgCasNgzUUCOhtgyQ35CxHiak3/SfZeCIYTZUyQXM
dr2IbuVCDbv0BlEq6QChawuBdZiFBsCpJ2WO41c1D/g+zPLiOx/4qiOuHXRe05/e
2+81ld18s8HQp7VvjsTkN6xyqVJfJe7h3XwDrWJnYbvaBJonqDGDNw5+oVqjoSek
efiDEW3BMfk0/0jFl3dwb3ekbv0vt288aeOp3iyLReLv/mrzejRaFsLvIE6TqpXX
KQnF0od+kNoVItww0FiwY4U1zwUoVUfpD4NkF0dKSWAKQCsNfeK547aKDUd8U2Lt
dnu3PBW6wUfyIFo3kmQUXIkMHQ7uipr3iQPCC72HUy2wxH07j1I17ibJqZvQqwHm
kitIX0ofHzOVd1bJpYtQUc3kzTKYQlYg4Ab+FbDJdTmcMlupW1nXfJ0jJANuZp2j
McgMlhO7aOzrKuTfw3E/kMI1ole6BkqhWJpiry/rJw2PrZcFvnSiI5O7HwRRHdUW
LL78OU3fFeZo9IAZs07RyWrf5sriVm883b5kBbw+XIgtZFdPZT67Gb8joOzTWSXn
ZBYH3n/FAhBB+/PW7fJj5AKf2YZ8IPIyuoskLmgADTqB+euf43LmFgu6Fe3iz70s
iO0RSL6N8SOLy00Qc8DJHMof3m0vzlY0Zt/mm9gT55G2UDV4gMJ8o6xP7p4yizol
Xo5dtJmJ4mG+N/X/lFdCSrLgGpPzc/FR0nChWLn1HyBuA40to7D+4kCG/eXO3tH2
9rfEs8FsY8h/+xV8dtPGkOlPJbLW8J95XmVcsnmjkXu12DG4gBU8/YLevInhhil3
hJBmBjPvCjq1eUWCu1QcvzhCrZDEY4XBvBSroE03XgK7vfugfjTorxKY8LixWpNB
zSzPzvmyvccrsH/e01/6+I1exT7XnzC2e6lSTGsH15cujNFdi+FKvOcWRSUcWMso
t1SxtJlWbYDSeCslDwcD70CGVS88jnglpsq2+qCxWqKlMgs0rwgiNoqPmId1qEEV
86hwH5q0uRGP01+VWtQZj88RvOxw5Iv1frvF2RxnhARR9CANosVo1CjJoEc/Epgw
0Q9CG5btx50W+SF/reWaw9Wd0fQz5IkouZczc2DOOcDB6vS+9DOCmsXnk4lw9fRJ
yvccY9bwTxe3qEdS2J5PHXl6kxoJqc+4ctk4qJcxcI2woCyGLNl1vjXwVfpN/yL1
OTLsoBHly/uNev4F7Myc1XUqXH7gu6RxIJgXWp27m1aO38rbvKwnpBS/OyzhYMtY
4C/g0u1qBBOiJTj/y2yzrZlyU0A1CNYoiyyfMT6kar32DR0TQDOKfvjPwUHOfUyU
WfoxCSZv8MgiK3rVw6CMTBf2v1XH+w+yksLEIG83e6pY9WUmyk83ZMDzsnnpftEW
9Y0D/9SJHlUE4UrfoN+nvcu4KctxX51Wwvjj232o0wZkwJXCKh1SEwZ1iQh4KjvH
5rEQPOr2PLlNQ4oLziPUBSKdbPLuC8WpcI8wKzFM4VFbDdLqIJ8wpQd6LRC4ZIQO
UxAD3KZeJUqaHXkeCoD8BP6JlPOazp6DfXJSjZpY2lm6RcStuV9O2cpPplmKLQba
rd/vDVQMYKUhvMQerjymPdCD3C5CSZTrWSB6RJl89mZuFuZKO7HiDXo3Tc5VslxX
av7aSkfXmuc80ADhd/J5iCUIX4E/3W6XyNYqHSWeYRL34Q9eOaIHY2oaQcGzUhjv
oX2ONHz/clBs+7aI/AOy+f+cSd9BpeWMd9Ewr9yEeQtwSXThaWnu6KBZ1yAsVPwi
8iv64y3fYRYgGFHjt+LPS096D6CF52I65bniquliPOTP7gCUfw7WdgmuiFP9xDMg
cBq1vOLAtcyHNP4fbH5mUILkgSr3W5G598JDyAz/BTGhBbV2ke2yoFLLyux/Z/ci
/79JVV9jXSW1tgMh0s8g/hspXpivacrGlfUuJcRwSTDcHtt5hoiVYXzba6/EpxfV
uHxfEwXsA7tsmOxpjryGypeji6C2Vp+s35BeQQKMv7rRaNRnNBLmZJsHgNqFiQfA
iK+uAoRONrAcSSJdJwKRga91Vea1e15ATF2OdOJxxDpxhVoOIvFP6hRXVBYGFSzS
vpVK562OTXw7LLBOPFJ9ELK2YD9/6OtAi68ePZ4XBm+gHu5PQyi5ZfAtLMfE5qhQ
usdX6QXbKG0fPzCqwQcK6Hi5P2n3ZIzGl5MB/kUZb/kX5bXLwYXcUEkMzG/oPp7b
Tv769w6zFO8erttBFKj/K7xr4NkIJRFJYWZlZeMeleJ0OXQZHR6BAzpQZA/VGU63
496js39xkqAceF278NPfrgxeXIgLXsIVtadJ/3qK+KZeK9M8pJn7xWYfb3sdxw/l
r4RylmukydKvyIRf5dMWeFWm55U/iAhBHSgoS+vdH103g973QHazfGmnA+zsurQ8
N1VifdG9OWvzJC4D5fsHIhXKYBnav9umgnPH2VcZa9H2FMF9HnS/OYfaB/SaEdDI
hfghoULUjulIyiXurwAWJARqHktzdTWlb4FZNAIbpLHtVnoNKP69KVbDIXTtbBwp
aLQ9MFspNOSIX+LDOvwhvr/KbxrNFLIheRFq0FjQL8FXfG6RIpJSnXozvY7PFgJW
/a4Xo5XqkJHWBmDlgwCnPjPC7FQ0iDt7J2FMq07YsH3J+99OEVwTYge9inO7IPq0
q/X7Y6hNP3QcHGJHRsb0WtZoTpW3iIRDsrU6bkuQUGfDzVqf6OcCFwCzxxNBOio2
thBxHZAgZe88FPwIhiXMs2jlIBUFoTrQqn6NPPkRjkX2VgNbtKwFKBVktG0q4vcx
0Sat8knyzfajqWkcucgE9aP9MppyUo2mdbf7G9TAJQuPSaF4g49pQjtnDKJpEuLm
DFQlvdgNiHwJDzWXOJwEHPnj934lZL/BaEe5uBVsJnhIO4lrqQBKweSx6ixy+b5Y
4hiBhY8oJoLZ1PyMqGhfUu6onLiBCnJOmpkqt8x5Xuf9c/+KEFiO7/Ictkennu0u
QNe4P8DqnpC0cVlXea6jdD56D0FdD3v7UfqMEP6ARPwd/3tBM99YLbavqJFY+88P
vmkyNPw/L37xM6I8bekCOdZUg24BpygBx0Yo7T9F/bBgjN4eEXOsURWzYjiO99UX
8sY6r/xTIy5iOCBPwb3Hh3f2JcgTJOBCycPfqtsCw1fBuUO+CB2FRiB/yZ6zuksm
IMXB1bf1w6Mq0/H/H2CcVfm32JlqFHhSRBpDgI93HkF83GfpH7JuJ4xWqkVFW8VV
sTwtFzizYnVYdT3Z1NQlcJAsxBjnSUCOGW8Ob1BD1x3X+JOoLgvthiyQls/TunCQ
2mKJVs5Puo2IK5NVuCk9AapdfTWBNpjLMTnMrGIs/+svvbVrvY50y1s/d+Ittt/o
4HvHQeF5sKHexwehQnMXyjAWEcS3BVpgcNBxz5eEqHBcmwSzqnX9Y5Cci2PjgQIz
KhVNW/kUB7Bp2pZAR6jJZoNh94cDcURSSSuoRz/6t/NXyVZEyRUFzyMkGkkDfr/Y
suStc2M8YrWwz1KDwTCp6fyKnARTYJZazGbq2egm9N1lI74uz+JOdtH96npVTMc9
89+lorUa85VOW/pgL7/LFBuVvZsBFq8QBYEEWz0jcUKfMo+pG4944KoeCpYplpm3
iizTZyWueAkkZ3F7/qmKfROJj+FuSj7WLpBaK7guzWKPNjRQjvJrAWe+sV1U5wE8
epCRWSqKSsaRmpv8j/V39QqYf1HOD4iFjrQ8CJ8GU/lleowiCTOwMMbUehg2ABcO
a4lcILVcPGEnNOIQJiSBcA5dD+E/DGKjbsIieOAuSyZqnR2IgMKSDtBUA1jkw+Z8
5RtUKqMNjlor3rL0xGLWfs9EfMDBBi+n1K2hc5U5TsPfZXtePRd1Nrxn6oAiBL3B
V5zrLQhm17VEajVzqkomJts/ntUO4y7r7t/FeYF+PwJ44zLvg1aIFt5NqoCKJgo3
xTemlnItY1o5DrZTHTGz+linl0ohvf3+a02sjrKX1132ZtI5CUyRLpFdF5Ly5uo4
5obO9X9p9wfT6l8NnMxgKKbNeEzkr2aX2cKl8u+Xx53fCvBZsMCt8TOV9v9LGfXJ
urGduBlpE5GYidvrj3rYIroyEYWiOzsAiHFa0/MaYtURtYPXZd7MKjW7QCml5lkJ
cpFT1cvCwztPtLsIGSDXr8sdUz2L1bTj4O7pdVRZ8pH9U3xNMP1fjaGThfC3uEwg
G0Q93sIkjZF9XmDz7HsdDA0vsUfxv3oZF2YhY9u0QO1eD5xxTkROHYmYs3plGi7u
XPamv2ewW5c2vsw4r5AFnF3uuXInAHcCTbS2KvES52ajQXiTfFMQAKZEAzNBJRis
S4f0JR6gLy0PdryyAckO7wD4Cn83WidGMqjF+piMrhJVkXy6e8gU6xrIk5qM2eA0
fZfNrkFnzu/96KQrYaY7j52116Zj5EfPqKzg3ZGXeYAMjmaCHFhxeXuWvX38mBdl
S1j3jW8ChQ6OflH91S84P2cZdhNPBBdsWNiooh/MsR0o8uW2NmKHxwSsqKNDl65u
yHBnrCQMcpjMNc5GwrszSAFq/ebC2xVokAcNiRXsG/0rknieqbxrC00txetPXsEA
FsRY+nndyFdyvrA9P4vhh+BIyVWhMWZOl7hd6Hzm3WcFyNYCAVrN7RkB4bSKHWCc
RdopexdgWbxpRr8xUfkWGsH+HMmjXPkjaQUx89TJZaiR/XrW1Zv1t9FvooTcWf9/
OfhH0dPPFUvXx4+O2TIoVN5BBTsmMFP6AS2VPG0ecfFfrnmXiRg6oBiRH1DkUMG4
4j0JzDYFo92Y93NR4yS/vkJLcAFYTbNzPV4xhcI5Fuz4M7dq/JrierLp7YboKgmd
DVo400b7ir11TzDKJEF6z/LhMy4v6DLP5Q1IediIta3dlFV0QhOefc1ueHl+aDDI
WkREwboER7AxCuNW1x7ww7y0H+iA5l9SSuKwMTx3J5+FiZlBIJBZY7kEljpLEVnh
gLHkpqdhQnk57ZvYu4JIxzBIyuwJKuhnd5vFrkOuA3bbRk1q9r7RGSCoUFXNLOhx
dF0tLHWQOOnRUJVc/VJcUvFeO9GMmatqrevugk/Udw5UJ5EzTwnwPVEYOIXQwLai
x+uXVIENa5StFbAnNkCyXslK+3rA6op14KLKBBgc/02f8/Vm76LB4q1czlSr8A45
UusMwlZWnb0e84DpIWHfL31y57PGwz34di2e7D2WSLJNPpJDfhc6o9xZ97QbbhGm
uM1KCN3VJYYNN8CRm4chUGe1K3IHCBQRiQi7Ea6CN/Sb6PKWtW/oK/61ZBG8AvvH
wqmC2VwjrdmsZGZzH1z0v1xvDvfLO6azC9Y5lf3QbvgY3xEwEld3UyEzi44+gooK
zrXnwJaNYEKlOkAgokHV8y2YuDESCf8jvt6nSW+5t1geppJ8yKhtKRJwFVflDFDS
m6VJ3gz88YubZC3qx1LZ9TDlATzn+6j9I/9MHFhN28Wk4oQ7ISsrrc+9BhgkE304
o1g8TKKHzRdOnGSL/nzBGB/IjUecO6ixvdME/5t+jeqSWDkpbwvNGp7n+AaCr3H/
AOP/Q4cdSwtTCrJU2MJB0J3KC3cnILfNXmB14mwXl8MVXKfUQ7p0ryZTy5+ksEgR
VTSBTtSXLTF6H7p2JhNu7/szL5hSjOsgXH8HfVmNYhbe4KmtnepA9Rddbm5G1MoI
xoCANoVHkR0iCi75rt01JAWSn/N/UbUzkk/2atrBU8jWw/XPBqFH33L8xPpQ5BXV
Lcic2N9FDau/lPzV52GnWs18Q0RcNJFzIZ6/iCco+UF2U9fIfu17YHkub0eOO4o8
Rxe9BIyc+Cnx/cJK92a6aCbnDEIeClTB3S8maIYgPNVv4/XsE91Xjv0DsKGmZXVB
D137nSJlQXfNfzlKjbgAEw6cDFRvTbWe+upLbL6GlcBzqH8bhK9oNNXIyRW7zPH9
a/d75/OYk38WAkRff/f3eGPzBm+N0vFVTUnFk3PYTK5X+9EDKyZjQvv8KmY1ojT1
TT40n/IrT0HC4rvLv+vz2YIZ0SwKLzmrQVQd+roy1VgBUpWuVXpGDcqB4yPwFiLK
jZzNyVPceMJqt+31d74KdB0z4j/o75tr4LqsZmX9gFSP2RZHZPx4uWA8STJ0Au7V
tONpv99LPLgd1BEEPtfyIao/3koNWx4D1lAzQ3EqWN9QGzTTLB1BmbucW60kL/n4
x4QvQBKXMt4HN7KWBMRJOKNpg8EB2IGPeY00UIzGVMTKs42TTYM8i/SkE9uWGEcb
RhOOr3R52zsvkD5nm3fo8uw3YImLDyBMQTS0aW8ssw3aoqzTKDzkhQkg0YAMS3Xr
DO0GFv1kId2KLiveh3npI9pCgKBhEKLt8uto5l/KtojE/JaAHvq48Qyo8v1pkRpc
AuniiTFTddZO8ZrRbzYNmUDx+hQs8sz++UvsEGcMDNei6H9ooC9EDKpRafpnkp90
xTo+JngdMTDE+fgka2AhljaiRZn1HE+pzi7HomJuDKFQJrnz9q60GIZeFtMgphUe
GlS9MnQYqzNMyztafAJYQdSIFBHwbTqNCjnvrXMhbA2ocXPa8ra2jkiV4+3gnRb4
waotuTE0nyAcfxWD6+tZ5DXaiVV2Ac4xjcSg6ts+VjC8sSCO8VVn/p/+VvodOohS
SMjSesDuviQWmEAoZXkWoOiJFqlHtppxQBVSqXPjuWrivNgiJGzOBWxtqHUUnxjQ
Ydl1xrWsPTol/uuu+wR7f17iwHhA88ZrxkfV8A74NpNaNBVay8LF5+Ij7TGWLpMm
Daz40g29NuXj0J+wxdQH8aR5sjIc3CrVvV+ZyBKbUG+HdRPRNvriMuNIK0SeQWkD
77S82vwP9vNhgHqPCkApbFgjMz7QE39wqlLPfMNm8sfbgzHrH2bFdssLawvufPI1
3q1vIqVq/edmi87glCFXuz7BMqB4s3jSHU5aauOUP/zygLBBIAn73qPCFunaKCgL
K9eYpqfow+wY3xeOvwJrJKAj+chKZ8DbPfjah6Gq7bCaklA6Aw2cPEJRQxx6RTNO
FkEnhIp3Nxcb1jH1z3JgOhTNiJQWgJuznu2H49P1qmmkF8YSrq4Xf4Zmh3yX+b/r
vk8gjauWMve2sbv+qudiavL/CP678EVfpWASa1rU/I7ovNZWhzadZ9+2GWyLvYmd
fBErrjkzHTNQPW6zNPfZ/23YHpwr9NbeDhC4DeU5o3II/KkARHa0IOJi/T9jIPfN
OWot5vEJ8NR8LWAH/Ij0Eptnd48TA5bgVgcfTKRvnfc6qD7fgEBVnUxAyNkKbgVO
ft4Odmy+dTd5PIL0e3AMrqcCFqxfUA2pdoTlxvJTcxXxvyqNBlWsXs4VVJLIct0s
jBVEL/OOByz4UA2UO10QkHuk/tK7TsUlDuCw/p3dt6gFQ5iu1CghWwtz9cmvcl1E
+K/ZCHijjZP4+i7rLounrwT/R1KTfqM5miPOioX+KtwBWL0kSA1svAlMydUjnKwD
ERTktv1Bf4Xe5WweXrgDcJ6KWPBOr5gJmDqO6QVwxDN48m2OEp3MrnmxZHYYvFOx
lNmgt1qd9TLaWCZ5hE8bxll3GwUsZvKdbtVSnMYP5DFwgDBZqBdE7vDVfVRjkAZK
ql4KnVFtOyDt9SktieniI5+xRONXPC+K08e/MLslTBbHwG6tzo0fYZv7CRGMxQzT
KSrxXuTZNoCJEzCtHw+ngHc1QfTdDAXDWVi639glZftk7hPvdkcMVfkIbTegPowf
9wZdERrCfdt7Non3ee5uehzVrVtxwNVuIpdR67omdG4EkI1wjXN2VC8f06qP72Qt
wGVJcL57yPIAJTsOS7HCd7MxzDrMJpoFRQ+bXirw1/KDCYkN0db1wVDEXXYB6M/L
rjSzYTkh9pvDzEkXm7wmXE+a2KdlqXgQ+uqKHiqaD3tB6zGNDxgNMWt/PX+Wn6cv
KAa4/EMVXXCkl9c1h20MkLHMjEmESY4fagxeOfUfo1sMdGFDrO06uFI7srnn9XZS
qGObGbDdKqs6G806kzX12szt7WMvDqgjpZ2BbQD7pFgZllgtkcFa/j/yq2G2Jy7P
/+IrKGkplw2Ke3pHXl3Dq/8G434DlPkP20Zk41HoxYE8rRGsEMtVCuXpInMAbF1r
gIHrOUylyR0KQ0ToU2b1vvqF1WkzvRaqehdqZiCSgjAezmvffbcSYqNP0qQ5PHyP
StsoIKw48dn4ELPkLHGv4Wz7ndqvrF7DMI+qaNVXtEwHgVkrgau0ddyZ/HKtGRgB
xs/s/kOrV0jrnYimJH6T6QEmi7zS/QCfaTXM1w5rTm0vx0qA9Iy/uWpLDcSMmngM
xJRMPceWttr9FA0PpY4q7O/3jfU1/HmUrGrWEhqDPfK1ShVrgYvO8oq39OzXm84p
TAABxhZGUAtr+PCAL0QiMO6xBd9S+Y82NwG3dmdSOqP68no00lgPYmiIWvv0UICV
H306XFJ2jzlTOyg7+lhkfRgLn2hhSvgvPE5p456OClgIwhxIRM6g6kKNtMVXXMMW
WwSc+ioE0O7XXOKaPGXZ/YTQUyn2LTiL1HLMbt2Dzn9bE0Y9nuAlj7ahYeVHtoOS
gFiv+Ycc/WVhrdNmjzYuiUZyoxzA6bqEzxwMbO37tfVaNbXcnxql5eTua89Vo5Qp
opELHE5rhUDkHPXGF6barRxLqADl0iwdtuRMj74mWb/4PX4m5TxVOV8NAB4ZwWTF
vcZOHcAaxK+DVCAWK5fnZ2+6qY1y9G/nLdL/4bACiWE4RJROiQdi/ZUY/SwnSMQv
MQm7y41coOdWKdRbIEh/PyyDYoJeGbARRxwhoJlc7xBOW6akP60iETKkv78zDurs
4BiIaCZCMFMru4q34GY4Ld5S/QKziUSvOtM217cSI4Aiw5LBwxvuScWu4ExbSrAt
/qT64WBibVr2MTqUTmPrH5UsrWwbH8nHdM67WNOkkru4tKPGDV9ZdqOQYJtgujB5
MuNM4VRs2iR8p3nNl6EeyBNcAdxvEvJbw1A2jau6nTsEMam/HqbELnOxR+tcJTcV
ZNiKBlh92XDw/khj5d3LFN2GxXugWwgpDWKBOaP4b67hyq4FqJwVSJyqR9C1E3vs
a9sys9KzD0a255pzOkAp4Ju29dAO3c/NT4k8pB5NEfmoeTUv6enDc6vPuKEkMlnN
Z4ZyeLlbUo56asXfR9NjBIkUF/0fgEn2Q+dMsyU6aOCebAzKWOJEyxgtLzO6RzfR
VkeOuYo99Yd30wSH05Rohm4Qf95+0blpo6VVNhjQAElruDWcMd7Ywvgs7nSglbZP
kQd7ckdrin4KJlVpbiCHmQNz5JbJZrm+3NY74q7nH/j3aVGcna84NYbgDQFOgQbP
WNDY0gVZnmyV7FVfcsNJfkpL8Y5zCzJWVJFbspCJ2NMo8iDOKKITCAUIBFxK4loB
uHwm2s5K5oRNa2dcRcYXQX1j2cOdxLe7m1cg5/O/oNAu3TxpG3JYol0xTsvJlUin
brephhP+cMPRrXEQ8USVVBMUXb1OIFULkIQkizSZiAjZ1Q65L8xQhZvoTwz/gt8J
1sNBCT3iyE7r0AY3B2VwkAWQ4RjZY02KH/MqiOp3ZpjraJl7E5O3lYuVrUHxohI4
AT/rT0NzDH4B6sitXl4dFxmdJGk7MjMbLbmKhuZLC/sOxuRmyiESqmwQu3Ztdu5L
tK9PnYaGONF3tQTpxYpuL0iqwWPBgpDefoL7NtrWwjz+r9JniLHp1y1aHGU0bGY9
hfya4B+KYM1YjsVIxqfKfdgsJuhXmIsW3frsMrGBApBh7TC2dI2rPHy8SztyBo0D
vuYVO/r9vBJmhQsb0+V+uR11EC/uUZrbDJj8ARgJNzWyT/S4g32+K5PzIHvsed2w
jq1kvpAymHVeo174zNexq6r/HHmnHC5veitEAGQs32E4U6yT+9nFM6ENCotqsmW6
cvTwDzxLoOLti4UsVwAewl7su3K9dZZZSZRBpv1fLhh/00Pxt4js5e5EDD1sXwPC
xekDZmQ9FPlJqCsE51DlQBx/7Gz8m5xMGzC/ifmwMkuXWrq1cqvfh4DuU5Y99FLQ
V0DEF2SQPUw9KdruxYl7t9YI0pI7xuJlJux7A79cwFnp/EQZ0Fq/Csux5lyXNm2C
4LiGiaJRPgjfOcW/sZRMxQp0t/GRJnS4CLNZEnUmga+KBVCV4Lt/a1uymi4Mybu6
MLid6vKPYjNeK122LXLzAf2Unr4RT4nYndptWgmy1/4cb2eiGbnM3J0cvff4j9Fy
hDTVLGeLktE/1StWNoHW7ej7Bo7PurWQdaIFGB7Mp+McBVD9SqvKYxQ8w8bXg5+Z
erxR8zZ4MArUPGHySJxfMvSX8OuT01Ch78ryPzJdxnq+Qe9Gm/Zu6bApjSj3EeOx
z9rklDlBvk1IbNtMU6GDenkyxlmfcj4BKf1+Mo/6LuiA05E+9hVjQDKLat5Qrc6c
lD4ypA0DiZerwoY3egGkQYmxk8x2PHVoZTa1rMTqE8NZHDWWFUM7+z447JXsgLGU
0fgL3b5xrXEjhgJV4piETH016opNWpF35VQ88WYNIJlXBuW641dvhMLelD+qYGUe
C6WJud8VpLHA/8gCt/hufx7Xy9Nq11mpWDrkGt5vGfGG2BVA7BQxjWcuRFoVRX86
H2txcWGgR2ZiABZ8rHtU2n6IWOak1j4azqEAv72GXjx9MYa/qTIeSvyiWSmRl/ut
VU7bOy3DQvhGjXkZ+afxe6Gy7xAwUox2ULxtsp5j3iILBIuhtf9dl3Kybz5GByoG
+MP3SBJNGdXvEH8TTHkd8xwtDEitq7tUf8ALP+ShLvBNAHWg+A89oBQ/RAIqIYHy
o2rQNHwL+sFxWr3h9KlSRfmXYTZIvieFIOtEgbzPX76KADZGi8jkX87OEzA3vqqj
86hRbR8Do6eSFn0fwh84cjN5XMD7Lua5AVgUTP4pbbTTETGu2JUvXGMY8tFx22uQ
GAnZDtWhD3ngNgpQspJaRqkIVYbIcAGTWYTHRxyVTxAJEhFD6U+VCX6YVWsvn7Gr
UM3NUXD1gjtfjrMbByMIK32XuNnZaOB4BTs9a1Cm3WqMQLmwD/nDWldR9NTbCMr8
9J14ieqUQs/o/gxxSiQBmrqrd4WFHl2J8McILXP0NjJ4lUxHUs6fuIvCmIyyzkJL
xOZDr9S0zOAgV0dYtlS1kRBkCs6A2jwrx3gXYfwjCqB050iSpEM3IyS2ZYGtsOE+
+oEkjZmfmqt7tFe4jGEgrtQ5wRjhK26iajNhG+f1108pLidFACdEdJvY8ZntSYHE
e0GGJlOf1ytUB9y6jqkeAZdElluKsNv3e/Oid764HFO7Y3SXjYRzie5vIYIw+ciX
MtEeJF+Y6z02uPayvABgRe0RrpVakiMGf0Q636wawddkuyCu9pSr77HMMXK4iHZF
49dl9GPR+DkbbRRlDz/qY0agTPX3LKHda5HoBc3cEPgx+QwXIVzAjKFDElt7fFgu
w+QTM5Ld3Fdp9T6gyixn+PsyPpRiDn/88GFSxI+JPXBKCXFaYvLHdyusRjsKpwpU
tSRctISqS+uakM2PAfP0nQBQNj8oR22BQswKooCpBjJibLXPDnCW6QcSFv/VJ7K/
R3jx8R/vORUKah5gs41iBIPRBYN7RlKsPeOJtlGHy9XWaIhqP16INbnud+hSog4w
5S1t/Y2ZcvuEcHaC3Fw9nliaIjakkow951WGYrUHmtNILmM3H/51+LTJ17TgApxk
KdsWsRFtWmdBHAqnrtZ13Vm1lbqxM6+pAiQLjnBUkDDqYjQO0arzsYNbfRxvo/RJ
CvI9uvbg5j/g5U8eB0xS6kQ+eVXvAVzM4LaiK79xpdEpigVAhCfTiQ0m7nNw+hTN
pTyF/h1zoDKlqLcO2oHOf+pGJxLPzhlEl15t+P+/P9+9E5PKCppAcHtuHhYaa6us
wHIjf0Fdx0EeE+mr995Fsu+jCtjsHuXNNkdCrm71qPk1tl/ZJmmSbt4TzctNhIfp
B0McdhsKqmGFDTY+B31WK2dlEly+AikK5rYxtDgGJWGJHU59Xw66X8fZS04/SjU8
D/lLPJPRIK5wab0k82xp9JR9yf6fFx40b+3dhzkraJKuaGC0P0Np8X652m60Vgkq
3zQD05VXGFZ27pbt+3EEmKkR/Qz4MtiGc8cJyS8og530lVLQTd6S1wbBPGleQ5bG
WhmBwGSMPp9TYJAGH25EbVPKWBZK0WuwYXY5twCXZ/tCLLFNTHJ/OHkBWwPjun8q
8d14dp+CKqj931710ORNfHPQ62uG+v4G5oJAm1PDbgkLJYPwHPxgUt9itmN2se91
UJTKrbUC9DFN2QDCkvcNbSYdAavugOytgR7g2IgLmHmcnFkxtZYpx2FJp2OnmJyx
VU2eEjdjGic4WuC3Hs6oYWoABBIPgmVI7yN1U9vNFmoJ1RXVshYuYjrAYbjGtDjZ
unbq2kar4e2oGBTo3uYXEDpT6uPLPAhgFNEbeNzwHRRoFzuhdaafYFBuwZcMVqOE
/n3XNtzX8wwbArwO/NlJre2TfGVjE1v/h8Qehmfa6psO/zpARj3bDh9lr8ZzoGAv
0ZJ2NnDPuGcBg5O5u/V2b6C9VPcNHEhN9XAVywW5gRLeYzpayXDWCXQCBg4XHp0A
eeqiVAcUQTPJ2Zf2TfrrZMPURGvn8l7sZtelFsVhTkCsXKMp5e8sMGi81W3lh8NF
pVlKCEpTs3Zi8Sl3RrJqAVfKRehYlDa/ZUQ84T3BRG/IHfE2MTX/FoZRqoif/Avp
GI13NaYkpImMpVXZx1EG7MVqgZiICFC6aQCHQtYlqCADSDO7wJ1bTsEJbPz58tWQ
pGcpaTWxjbt1tOZfvmLz09jUBCLZoj+U216VLi6Mxksn4c8DcKB5g3T4KkXMl2A6
RHJriMwiBfcp07NgddO/HMkrUgUtkyhv/oar2a+l+7ESKneNJg590LCEVI6av32N
ROPXLuk33C1gqCeMDwoJKnsprKzQifxUdfz1xBwLHIqAkp5JAWSeZlEetP3Wiuro
Ca2pwqJAgbzgPzgEqH25CAoCY+pUiZq3cofw1VvY5BcaqDadm3KNcDKzSsHpq0+I
nVp7vWU4LFi9IkpZxoQ14Yj5O4GtbTLnI29mmRK2cnI6ma+LFaZ/S+JjfwIXTRFI
W0yCbXMUOJIEPT5HBwO1GqHmRl5tGDMiuMWsqM5h7LM9BgLD5NAkFXQujV1xsT5r
hJFwgaDJCB27U1yE/oFxROTlaNfApKzX4gxleVFullHrG9RYEFWGGaHZio5AfM6M
e0yAd2FG4v0HqhfVC2OhuWxTnx1pE679FySydBa5H3OatiqWoqbVdYP3ppqAwiAT
gDrXrPFxGs7hnblu1epW1mBB/2kwaMshmJDegq2rdzOp8AjsM2BMuxv6Z/C5RKoy
ZN6s9V74Gy9s1mfVhE4NtZHsGowFf2ZYnD31r2LWbLGo2UJY+INIk5oNo92UlThc
eecF/vh74PAtBxZd4mnUgzqvZFnQA1eVG3QQoxon1JguSUwpm6dpj6Kb0GTZqw5o
H8B//5ec/u3LIMyzZ7sWMdjnhYeyo3cXI1iS3pzZf5gqB3/Ti+ptHVLjffSNdlB7
6CBV9RHgxCVEtm/8S4j6jVMpP0NyjUWKXuVlUKrnbOR/IG9v+2Fh8RdEV1zcmouj
iEXzI8PrGDlvJtxGAULEO6Prp61qnXCe6yziyJFJbvs2+BheFB8QtlsJfqTJ00yr
I1oaIpW335T5ZjH9chz46oBy32CYRaXEkb4Jy8Tq4pZQvOuMrOKOgxCkIt41mxLQ
DKlF751xW8DGgksFAcEfF8UwCqk0cktoRjB2y+VC+u/q6K8xx9iQ1UqkmheVDvax
B5vJtkYNsO2s3U6j9sKY/sZBmG6TIh5XHYKJPGeX1wIsDBr8darPTdiLkdsVHJ+n
OccUwM+FfO3DnZYJ04ubAAPqVstv4nGUvjj+Ng5Cawj9woQCEACOrFq/syFT5jyP
Ijj/cEi4LboIMzO7IZJvNhHKSdKbPcs8VVAueG0DoFvsS2rM7H0jxoqiXZLAFOwL
DQ7EBWYAM71i1UM0CMlgL2GKmlgeU7OLGt5IjkrajWV+xUlfes2LMZsdwpA1e1Do
w7cH/QSaK1FWRU6ctaSSxS+Fa7HlfH58SykeFFpfa7P9Y9543aACeGRs9T6x8Tww
yJlJcaB+tUe3R7JfG/8dl5TgACGkuuZAEIXIURNVJmbzZuI0HE63h9VtSDVcvjGA
C4tEe/ox+k7/n5haZ0QN3MIK+YREG+fTNsWpxcXi57Eqgehph+TALrC8atoXnvlJ
aamZmnM1zv5i061X5z2MibuXC77o7yM96L02YFf0zwHfOczCFu3OP7RXH51Ld2yn
QTw/eYEYKHovVVBk2QO0BPzLIdAQEnGkx5PcwE8fs/mceEpaIxFfC7SDYfYKjetZ
dfEQdZuEapmuiB7kWiIb+1cqdlgRs/7i09JhucOAWkadsIhjBqTTKUCWYsEudLJ6
3PqMuFtf5lbCdME1NaRcTCRJxb9/qeqI6ZpMUOw1njV8aYrw8edvhdm2Act3qyMt
/NgRDvr1dL6qwzzJMG+2+uKn6qbZ/0PFwoxNGJfSL1sJY3K6kmJzo4c9RqSKOFj6
g97WeQMQLQfkg3krrixBhXpwxnO7We4UeysaT5NSH7YIHgj98kwalPnyo9Ff6oNq
KqeMV14l6raHbR7A6qwYY0ldN1A7ou0ZOrPP7PWPWC65diVdaGC5YphjSpvOrJj2
WHkjBMHGw3A3HL15HSH2LX0mMbzWyDVP/PvDLcqztIhmrMp6d73nMD/FmLIsKUN/
BGctW39zHavWXaKMgsl3J5HbsVskunvRYmBxSrwFIts9ukVre03RjTwyJvsF93XQ
0i89gdaJz63zsAwckhWc1FEeMWTHgx9futs57fKE/10LHzzQHAXDhXag6wtxbYDC
LobrohwWT41ZjXdo6wn/bb13rsSHG+gNRnY7ed+0iemNP6Sv962SZd/u54M/R2iZ
3wnyKbUNK9uyx7FiMTV2ehNWzUyLxX5bL8J0hAPRzLGMgkzoKALKS6S3+4+FwXkK
cT4qmAWKa75KTvRl4a4iY3qOsFC6dOuKf3yfAfICkm0RM4y33I5cRSrSHueebnv0
Q5qshslPv6qQFfmdu2f3Z0qhmADJSFae8Pww9tCc/GIZkBWNaPwaHUHQnfYU6a32
LUnDCJiHBJg/FhIJxL+OOGtHqz2/rkEiRmnWDN8Q1U6mKRj0D4+sP94/JcEg7Ua3
u6605/1AM1k5TIOkAqaiefULzfOC/cjUa1thcZdVF+QaMgOYvpoFkIe0yxOK9F+L
j2gObu6PUIK17+6wT29ks8elclmaD3WQGZp71X+qIm895nZPgJx7/YQwQ3jX+qS1
FxiL1jOExyKu+JkYgubeD5cu3wMae4/1OOL1eK9UZ1ykHG5tpl5Af2879cgmkJMM
Zjv73BL4SFrwZ3s4+0vF0r7ixU2EGjeuhuFxAHdqXAceB25GxXqfqCnLduHRACZk
ukUCVAr4l7x1QdOQUuL90oK1in/sgQVQYmG7rBgcEaB8o45MCbu57d5kc5Wktwod
t/NGop5Lxqw9QBNfU3HlSfzQX2ALwi66UwR4pjyhZXB6VRa0BsdzlS4V/oWIeDyC
zW8AP60jrxDNTz705seNOvGDNoLbNxRhXhYilvVs/Uyl9GOJAfofJFExjgjNGQxw
DHQpigC1u2P6rwrR22/b4OM3jK5s+6DxLPaFf9F1GwA+syq4+/0dUiw49pitmPlw
BHYeXzL8gXrMuzUGrJgYYhqm1dUGhXDzHawp9G/2cDYzbk0I9/cRohEYEaNABs2M
8bdKb9TPPJGqYt3sI8TxbWggXxBOC22EQXffUh065ZeHZ0M8laXg5unrB/iq4olF
9WiqyUPMj5lQJUAFGT/3fnDiy9Ah7x9OJP0+AiU3DVn3+F3NDwoeKu6wT1qtxxyl
W507LKkZrzKhsl2SqIFE66J4frvojYw+V+L62hWaGJbbmlDSuGqPlqAR4Qsb/7X2
r2L7yjsPJSRU0WbvTW9rXSkfROGo5RZ31VCWO4UigjyCQtE73RWplrNQtDJoXA/0
xfkXwUs8sINOhU7ytdXqm2OvWsvEU2wmAjHh6SYz+ZVlejh/PkyQlkpvBtk649qb
UCgCW3D0Z8AU5imhJZE++Gamr1HEwEQcYuHuBXzfExxiYph1/Iltwv5xZc3pybLB
xyRy8BNIKmurjsaiW1a62siGqI8yG/1rozJPpvHklZKsU7iKll57k0FqOuZ7Cy9e
Ygvr8xlt5S/SkIx9McNW9UTYezxDDTl1lOiHA+yGp1b6VnpEZLv7Nnq9QxE/i3r1
RZk8X4DAaTfBilDk7UNFPsH7n3EMpN4mfETX3frJjKSQD9qOMd8jStZOofGhNfIj
Sw9e7erFC3gU7rjwMl6pDGtmBFQvJwNmaXsg4XUcSQCvLZEyK21Cq85ARNX5G2bm
YndzxkDUY+gm4Zx9FN4lsKZjlcQ/AtwPVA602MmuozAnxiTJ0KbTuCBLxyFeF7Sd
q6rlr1Z6C+uWoE1EZB8Y0q1QG43tQFGJ8P+F9ndeUqIGx/RKIHSrLYNFd1lhx7CS
R92qaikU9Ehwm/DJv6gTbig/pF/PQnS1UOE3yafAL0E1dJooJ7xzaKSqONB2AsUn
Q3lih3KIloUlLAsshD06zi9QbpK9KBvQJsie9slCKmzxOvVYl7nDKWzUE5mouFdW
F1YI1nsBWVJQnUodNYNDdvSQXbeWZxqcS9dVhfseJTC9S1Oab9b9SjiT+LFhYVEs
mZk0KOHN7+zOA/af7iC57YWv+XXqCCbl+CFp7+v8kwd3cwVpztiJ7vEpwlMW6mvp
c6Zj5DSy0OXMSipU4veI6ZJjIWTr5XswM1qZ7dEL4tx2zqxqlO1n7R/IyrRnXQqf
f6x/v7vnxEedIXykGA5fIHMy4dF16OHR3RSYFB7CfPJufrXcLnRAdtrRL7Q3Q5dH
DRZ+5qYw2LMxipzRTjp5OMDu3Khdy3yQWN2qmaKvd21G7p6FyfT/caEOEa1Ymc1c
wfUWcG9vYJvOtgnlA52Hu6mwoSWro2I+OhHURtquItcEhliZ+gxRXwDlPYY87zp8
7DBK/B+ZVRobgQmwOOsVRz0tan/A8Xq6TPwI/i1r6M9uTTBe0NCnxunzDkjzLOVc
ZhmqRcglM8Jsyve6UDFbzykaFRkIKVTW01NYUgX7LR7FJ+p6YOzm1z3KcO2j1TXG
mmzz6w/lkVxfw2kNFvt5PGnp+/Hhq04ZqAAdMAGROM1AyxXsoq1Zbi0pJJ7qfChK
kJZRyWgqy3HrvZW8RP4T7heMK8Rtyzn65x60HGqABybYYZV014Z3+E3lnA3J5yZn
kwFt5Kq3hx8jOiJdriM5AIm20BFV/GejpzZkVKBGrntS3kDO+te1IZ3itYn9nA2W
TNwQ68fdvaATRLwfBXxjDce58upNMXyW9deds0V286hwdTvBBtXaTB90+OYn1uNl
PIDD/dDe+1+JRu3NXLycbCRuGYexgMa23HvAVKfISxCieK077IzKy/rVdV1x28JR
yDoHp8sQ8UEZ6WeyKQLnZTvtJ8ukkBkGW5mLYFyfyVCq8xja6HmBD6hr7mGygPQq
82Dl5/PlSb3s0gRKEYmUMRRIj0/bIqZYT1xMcZVt90B7fJIc/Pw3KBSdf7QyU8Dk
JV3qkzmHxFzGKi33E3Pa/uV/WMTnFhWvfv+/4UXwzJX+JZ4+YpWRxfBQZgHWt6lo
NVh3sKPpehtFEOKJvtyKoxNrkP5EnDphjEdSL0iasHscgXIp2uKy8TlUxby1w8iD
SzpDXO5MSA3DQ1Ydcc+VMhHDRgm8NnwCfBqifKPmbBlrn+3DtfBo28wUqkB/xAGQ
NLkGyEDcgg5RdyMqoQtclz5h5VvRKf8dlPAvDG3ik74DptYiZuGbekXEKAvR6Mu9
oowscbHD++5YULzrjb44EGbrKYwR9j+SGUGfl3d8jgFMtZvwwHyfqVDBasS7b4ZZ
LLlZaeZr3f8CF94rPX4z25Rr0EpcKKEM4P+N1jbqhwGMSV/rL1wP0BFZxBCj0fds
f82ykCOu7y6DZTB/YJ4SkI2/NB+kfU06eEyrMSi0HchtQjGUbLyQ+xk/717B4Xp+
BIVu+dWnK03/L1ylyDqPJkGcFPI9Laf7VrWdsb6eTmrL6P7cjmDTHOusE5GC7kDF
IoSAK5NmZDXIfHgbRA5FVbDKwKEvV3gFLx5K+4GmLOONjZMAceMW7IhE4pydN46B
CnMKAP0MlllFRhJK9ibLNnJ7et7o+A+UYJEBzQzAzPxvjvxvhMUG7k5ea6nmNwyc
ojZWR9POCIf9yk6sBqU5Nm5wN/X9jaoTwFfOY/JSTBWr8HQa2b1C1vmtoV1zVLnu
mwiWH+gaSZDQ2Qfi1oPhoEXNtnTsgzTeUivQuPS+Nqg4u/EPE8lNZJKxIK32yKKY
QeTtALKvIhc3Ae7D9AgsBhZu57e+O4n7069TBOkOrm7VSkzqODa/7iMpOGnJxnvf
ivkewkyqSg0fcoPChwzTUyMcpx8F4FQcCk16W9wBpLNoompY5AXxDpKAty4jzEqJ
IYkUrExbdzdtlcfmFie0R0BZSnYv7kZhht9ZZHAPcNwRK1y0TFYQeI5jZAY2Btns
DSNThgh9ocWREsHsB//pbAcIYbZceMKEdx7tpF9Lv16v6B7QsHTpNn5YuIc35v6M
alvvjOqphK/OBPNz7SzyYor7aP8CqNakyUBV0PmSV57N1DwuEQ/hCFdfvMagWRTb
BPIcaURN7TXTSZoVjBt4wbVtH+np962a9a02o/JVQ76t+U1/X9Pesjb3t3LLqYZC
GGpZmROrKvWEFVKel6j8akC5bTXMDA7FJbll962nP+4iyjnoAui0u0/gPIBTFDyr
LZMWK4+FRUIIcVS/uxMQJ1PfpJhUIdrsKA1pb8x60k4442T3dsOeewZhCuHomsmJ
vWfGrdqJyZAAjIuux8Q8/fZfZRfHMLYfLWpKcCbCQBPtBH3I6kt6CJAfKQxwQLKH
1CT5v7fK0Lkq49zPZP5V5iRPWXfmHpfxuXYR9IdeO94sNF/pxLlu0stUnbM2C3PB
GTAIKTfkvLAQVuXm9rhb0F1TPxLQYmFccJTnXlan3siSpjsUDPGauP02e/3Vg8Yf
K8q53C4B/J93cKLGTkjlri5Vj43t4xq7kgQvz7f3VGc3L/lPIMyH7pNXUFmYFzVl
kQWNfab1+V1NOs8dOuVlK09lxaKbQLNIaGc7lwYoVroULO+CVTtEltLNVG6yMiC9
mp4IgCDwqAa0NXeiUE8KQ0w9hx6GOOofFnfCpvaj5LTUd8Oo3MiUiu8UhwiPrFeW
d+Iy1DDEui4C5QVtsSJ9xaLbSPHFrK+3xKZxKyAhv3yLxPf+F3BhHIjCVXxHcg+9
EkAVYKxH63b+kC3bpCRsi2jv7K4SYrxQoyGQejzAILiSf0Ac9j5q5L3J5cwlq3Qb
LqnOKGZsHFq3TFq9vLF3RKJ33AcH3yzdkkRJPSxMjFKlFkuWscvITHiAuiiHhy2t
rAZN8f+1PZ3KzLcqsfqhQQ7uKxe/W5kcnBcPLeYgRTVhDf9gBkayIfn3yIPd7A1c
riUuRly5imAOCiJM4dSFmoQqPBCAojVr/peM2KcD3q7IG4RlXjOfJPbHn2uC7S6B
rLh4Vk688lWxDJsQ5AwFBvBVrdap8RHMD/JtPs7vG7Ue+Ajv0zaOI3ywZCwF212b
sOawijuv2aSqf7GGj1WrRDsbex1M91KLizlEJDbDYlD+rLdHeONQxx4LHwjIr/9e
Mt+lH27i5JjWeJ9K319g686E9xuhBofPJyj+Em7Yjqqa0LZ9tBKyq4FAOK0smjFF
YQpTV2SwxiAWCMScRaeiGvGWPcd7lp8+1vh3dDKxlLQn+qGSPUkMClR82GbiwXFw
DuKoGL4+GgEBK1t0LXyLgwNhOby0ZhcOcsicoAMGjEuxkw7jOM+yAqH0qbLJBOge
4Xv0GFbaIqDHWf8H/6I6FIk1OEDIjHwYI14TvOXhLg+tpYEQ76FquWaqBn3qNVcf
+nqt/hWojVmtEa/THTxe8pdjgi2izEFzHsQbTI9+0sSYSeJDbzj4zGEhot/FsXv+
WuNy0jWedUrnKOHRMlBsyQpkc/eOIm6IFWT5+jsMAYxEQdxppsFjNicyEX8EUZkQ
Hr+hsOHXfaEl+9IDSniZGQjOEUGfXFzo7Sz3Y/wCA7yNiInRiFNmRYCTsUWDfjzJ
YshNOmY4vlySEpNeC9k+hsjIeE7vascplPBsjYmqFmRFaA6Khu2TQ3txNn7XMCTg
IJtLMUHKI1l4RQmDBHK3SOJk8yaC+a0S4sQVfsnJ7GHVlyYcQm4kt9mKSlXZm4HV
2bB+Uyc0gJ4uIufdSbGe7XOVgxRd9Kvc8VX6Ix5h4OZmLKwJ1k+CtJF3ezMrQ/LF
uIujL7Nk1vy6kkVWxMYcIYN9i2SiVCTApiBidV7x1EKukJ1pRsEBe+ZaH3221QhP
KH30okmOxw6zTHN4KJec1x63eKKpIuunGH+2UOXDhKhDsd+sgY9zkCUDDUzPlgra
Q7bscJGKMexy4TD7AN35EojsTWecivdJ/4NcAST9AVEomTuHBAWyI9PUSsnujLJe
nigU8b4n3ijR8/uo5aoh0cSjaAo/YHi9A/XoRb992mfUDBEyrxxF8GXovS7nlCxK
Ki3KB7DrBskjZ1y9W6gFsbbQEfGj4p8CtWnpm3c9ns3kKgMmxPlHQlehi2Rdub1N
X/qdZO3YEG7+hyfpXTnWFab9JYEtNWVgL1IZ5DzsqTq44arhzyHJTP4d6MdH6XGW
uj95CP19p04MPEF1WD0LMt+0Fk2VmEs3m7bBaYRXivhtw0HlzL+X77Jb9gh5jOyc
UnoxTapkW1Ta74Ob4HuJ/WlWWAztei5+KJitDurKEgCGrUG9iXf0JIJ6+FfR/QSH
VK3PHBsSuWCe5cuosbPv4ZSrK+Y6kS9Pc6DXfW/aVKx24D3gR61gOZPmgfIa9igs
OH8oh75r1BGBH53wyFTFntNgVbNsG8wyMauW2d1hd2LWXi+ixRxVclTjceOoILnW
2P7O9lvD9/SErKEMGAQo7WFHkiHbBypLOocNAkInlWr2eckSMhnPDuwu7/XmmIvE
Bu3+iphVZYKrhxliuhiSp6tJ0nVJE110Od0XEjREWVVpPi4tSPOiW6MKwetFJ7sX
m+AyHFDIOpNnWOA4P3sQtETy+giV2IQ6nub1NF6kpQk3s+oNszKAh/LZcYytl4GL
kMSlT4S+sED6WydiEcOVGRuhLUyYiw6/AwhLfieiRSJGjTSRNgRG1f6gRxLAikcz
RGPnOy69gG4rK/5Hl72Iwo269FwKWouJLIJYDAmWBhkFa+pqV5kXpYQ/8VN1vsmP
/ri9aCdkDc7+bf1rXpHoRufgOD2IZSj5Zk5h040tMXI31RdbLT4LoQ/LRfLbdZAl
AjQFEHMA3EXsHj0JxvwhR5+6ByOXf3k4pjp4bPI3ePEzARSO8r279B3pYstR+7Av
OV0Wq6eWxHuLrDC8Xe7sNpvcxPOw0zfBb6mEeOI/IKQzYiDedyXpFiIDHxrokmQm
3xgqRXVg3w0+LWOBUZyDuUYFJHL9hb3tUC4z5Pw8RdXrzOEu0aPsHTSdOVK80QMd
bw+yRCFQN2nCQbFc8bc6eimxAoj5/2WwOH3Y4kPFzEHqolWZ46t+xXuq4bLpwiOh
uW2xL80Q/4YjKiDrqZgZb1HutezitAVc/RQlPtKBYp3i08Lf0s7T40zQqO26nBy5
FyVYgZ1fZLvWI1ebE7INN/BkoOUV6m32KJ2phcEo/6RSEP96jttSDG2UPOw+Al/Z
leLcQZ7dOyRQM2rq2U9pQCHXYExPyrT1JF5+cl5PArxwl9xenm4iBF09FTRx55Ss
lebsCgDcNiL+qZ7fnIS/4853Dpl4oUA4z4ZWU6+0xQWwAIhjvDoHZyD55seuEw4I
jych1GpPuIPy0IeZ5P956+2E5eazKSorkLr5rQlG/SZBbDkss7tq8MH27dlc4MBx
OIVfUF3/+QUSgAfAdLa+84q9WxZ5jL1/xqjXBYpH3KfMhEtJUYObrUjxNJAW/sUS
O+c+yHU2i5zA+KnYXG6ja576K42oDQYhpd/fWedLmQ4Ogq7CRoTqKCneFfHApIh1
ndLc9QibyEfxUdd39wja4XKc/+1s5B36NDwtKJErORzu+NjouFzFFWNY5kgccrLZ
cSN41mHzDvJApodPxFP3LNnthvN8Dbqp8sdsx8D1v8OH0w+FEtved7nKqDXYmLql
BQkDIAKrXm0LI829qfA6Y5w4q3actGZvpD6o0/O+acYIdApzgCm5Aai9+5YZ1dgl
xdAp/7p6tjMP8VRM0zV5+1iT4vHWij5V2scleasnRqcp9JMantc9q3cW+PVd7h4w
SEL5DXo9gSRkLPILAYYHO3XLxhha+V0lvTkciRJgwm0PNAODtLjRp2VpRcTOCjj1
48WfxJ4Huzb7FAK0rCNVSU+Em0hqq6wG/nnGFTqa0UzvC+oEEVQgv7xnimpZJlY3
Xk8kLfPcRMsTUOVUgqZodrPPIR/merT13R5jaA9UtOjZ/bJLb8Q/KidldF8RXPko
a1ZfjZRNY4D0iwAz4Ea4iY87r1RUl7lqmWNsNIAus4Gqn1bVzGRbafkIRrol+8LZ
XNIh/7atXXQOSkqyUGPqlcJzioew7Nz0Kp9LTmCVXjsFBjW8BsZVFn2t9lyVbwpj
skvMrZ0AxvDSUcaDGHtMlqo86BSEbN4dfrjnfq8OnfmGdH9xNcCgGYh+5XTb10dD
hUeTruW+1TiMeERBRpYq8+7p/xUgaddfTi8VK/v5nQAodi5oVrd3kgF3ImuFW6mi
zD0vLL1hlRRXJWs2w+zuhu0jU1Bu/Vl6Ylu/LBUNFqMCuj1FNZHQk75W+BFo8c9v
0KLaWu7ypVO323Ih/VQH/Fp51gjlkxNJbOtWyMFa3f8fAzet1mhg1trKKfn0oHa3
z5pkyRFg0Cy0O0A9xYPMSlB85WajAeJ0SaQ+/dJIwW1VwwGaTs1SK+5uExbw+NSe
qHG//FihxkAZiW4ATyOXO8dkqJK1v5d7nTo5wQk4IHf12kcvzsy96nAcZtG2d8fO
Al3594Y82YLH57HxnaXg647UvjiNTzF2gHCz39eoblSoHaKxuYG1hCG3aIvAMtwz
hGsi0PirjPPGVgLO/XXYAqG5Q/9j2vSVSOeVbObXuCKzfK+JIsq9Fs9LEnGJRtqE
eB0/5nqulKdSIK9oGIFj5T4JIsqGD1Ml2dNmrfjjCXuh0G5BXrQaEmEW4hmsZlMw
57qTYCiyTeYCv3BEJb8IDFahn9GkYVGsTPlAo1p3oYRk6Jpu72Z8edmGeVrHTH2H
9yofqak5HQzegHz76fIXcKxVuDIEfpUJf5gTvTBmChf763y6Rge6qoQ3V99zx0iX
ZSNFj0AyX+XCuU4cUFvWp2cSw9SEmb0ts73NHcbXg5bCzZpPOzdV7Ce1xhuEveKP
RNjvYzcUAIsk1xZHXrq8OThEqjf6+Gmd0kWCi2Drw0ZpiEzAq47Cvmq2OfI/CL4u
erdjOD2ee0XZCLj+zdWDye2rYOf4HTeCaYMaGotGjrZKkQyUuEe3zcPX0d4BmiEe
ZYuFNMLa+ERYE9QF3jqrvgftcoDZSNL2w4eLRdrY5n/S3ZXvizBh/Gt31kXJG9Ny
pINjpU6BKlyl0GtCtn3PeWOr3tBShm3eSCu5h08ojoPFXBP9D+BMdoEt4XNkNGW8
91HD65a1dyvkla4yFxUf9W8DlnB8OpQXz84lZPnUfhKm/qMOINnPCnuXqv2nyI0v
3uX+I2VdvopB1U5Wc42iPeSWdnmo9ppG+FEYFROraY+7PkccLiSAAFWJsXSbUSre
8dkpxBoBUot9wq5RAzEr/QUwYw0/zKSrJjADBxUQPKC83DaOR4NNqf9qjU+XWzTH
K3WKksIQAetmhyV0mLHp3Rr3jw1XHQAbYp/fdrZUMm8B3FK5HTr4tETrp7x5T1lT
I6VbUaPczJDmjyIl/WA3ewQ8KMgzSHhcmHnqo+84mXYS19FNUw086hY4S+FRNWFu
C5XuyLRTmydYQl6j/tM/uRSsBnppcjLXqrohToUQofv0or83Em7eI46zPI2A63Dy
ZCfKOnZa6KzDE2Uv8WrUZdn2/GV5E1uBMC1H2S7Mf77sp0+LrALGsUNv2HwfJIag
7HiGCAtuUK36jegAvxfpOOHi4eThnJuaDBA3i3MyFrIrNusMrxgGUvPCmpW43rGa
85CH9CBHS1BfX0i4oJvAXMm5mwIKz+mugtr+XE4cKJWG6N92+iyZIMxVV6995dVP
unLNud0vfdSYSpRkQyvnOlZvqgzh2OigQTYe8srwFNgju6Z4yIKtgwYzUZuZCjJF
JZkYt0vHNgzGn/xFYXlibaa4Klav5ejSlAXOJoLALmWpySTI2mvndl0iGX1FPeSL
FKA2UPGMDr68AyPreHTfjAG5ARu0D+2ow5EvH9//xY3lloviuKOai4OQUkpcJswR
8bmAMZpX1AFgH8VvB+Eb/fdDeHBM+L8qRHWJtT+YaYfFsDZGA6aY1M88jzYQLEr2
dmkeQKMmPDYr8I/SrMB+rIlvTkmB3eCmLgYNWqCQQvVxZ2DMsfwc/OLUc0ksKLbl
lUcYQzbZLeINHAbyV2J64PiCuuj8299vtAhJcWS1namqM/gbs/4dJ250yJje+HF5
XEky1/HNegDaoE24B8DDXT0sdasSqWDfLEKiyxzHpEEipgpsCM9B3PDfcrm5fI/V
iyt6CB1GSKr697Rn6QEB/jDp6QHKfVkLoxVg9FBjxjzMvZCPulxT4NMD49VjPej/
r0zUXjw46aLjjC35SO/VMSLBlTY7JPkU/Ue2bal/wkCi1t7wCjROjlEtdKQsIgz4
BHq/SSmdUIUFO6TX6VK3X2QHtEZ3IsEgVg2bt4plpZ/LDK0yJc8bAh5BizUSVMWy
Q6B1pES8KRgZKZWznIZfIwg/eF/A/UtRL0R1JaTYoLflTpTtcc7I8oisVKqg4N21
TwqqHWVpam+0iIySCwzSf+lVpqs7/oZP/WAndOgwsxLDrB6VEy3+VZeVducAhVT5
WKOrgc5AaWOiMSU9x3mAGM5uG0r2izAhT5l/JPn9391kwqoIGp9eq61JPpgPa1lM
dwxYZbc+/JZFwriVgwSUgYaFa/N08B3pYa0CgYQw1jMuisfGwA9eYUMSVNrENoDB
9rK8UhsV4H3aX8YEOy8KK62l5oy1LfOnsyy2Xztn0Qd3GApwbx9mEMth9Gw0SrZA
0BH0oSXAw8kqs5yvbOU9Rsg+9EZZoTZ8z90zSWHJfdjkLMlIQtJlM0cs4IEZmKGe
HwfvCHxy0rrmXUK92UTh/hjHOl8dxWVWM9sK11eTzdtYjTR3Ekj5PJg+u3NfpNSg
8jjYNts1nDZApoaiu3B5vHAUTjmUtaQqyDELie/BbH5iMBtZDoxwMeLbgtYxzLzG
Asa10Yv+usqc5oVIJtY4QzQGk0i/dVtewAu98UgyGI3zq3x+kcycfOekxHgXBRY5
6+UVs1URANSSTjwARkezwLrIvw3bPXa1T2vAt3xqzSF9hDak8Sv1z7tgjGihU1kX
rBv/Bc+r2YXP6+G82f2UtAcfchs6E3Z6mOR3wEWES5EdhCpU4Rk6zjP/YRQVHphf
ObGdSuJVSrQMRAoxong6p+4L8m3kGtKvzDx2LjCEUyYZpRB0LhIQPh6zsIjlfJ+M
PgjSX1FWAPI6gOYv7q91C6hVTVlWCwgMMb3p9ahuFnFIIwe0ncZqg5jiAtf6EYKy
K+L2UJbHnSvuV0BnFUPEaoI9p4QyyvBU+xjDaIhJsmOUCnbZNZXiC91H3N8t2GJE
YqF2MlpkaLyV/iC6p2c1UohyAQZT/AhYNjISIMP3kMmtdjXI1dvXfjpE13h4ZyRr
k9e2Ezt6iusdZGPzBQofRvPdi3myydf0w18ThkyzavGcEEnxILwFwaLpVz5/56fR
gINlQa/kd77sTt1gzYN7AD/uYHBo+/IfWlY5786lvYxpxRz44g/G0hs284Pj0731
BzNI2YGwZkAgcT6Tz7YRo0L2Vy1Rl1fqaO/exFr7I+PIUIFcHwmGOWipSmvCBpGm
Fkch+rlJRnRBjHv90tY7UMQ0f83Fo/eXscyxhAZktaV4/2LuMFFy9zMOufvyLUov
U+u6A3FIy1wR5qVFwyEniRjQKIDWxNDLydyXMe7LGMsx0pksR3QmijCGyQaYPiKV
yzZusxRM9dqh2URRqFZot9KKkXnAyduXniYWrt74xxyIcBOe6sMyYvsPRpz2bDUS
lJxSJt9FeGRAs37WN1PUrhuUjgK9P2k2I8YR5EjRWdtmOUHkbmGhuQUYuIgaUNCe
tdjA5sYbDzwz4VWn3XFWeP3h2PVfnGLI9MGFUljYrBlMmGCvQlglb/wBgqaWRoRe
PG4ps/XEN04AK/EKYC5zBORzR/Q2U0287aBGAizdGxPGnIWnAWPs7uUNxkIwOxG4
prwnnB5USieJLyMyZVU429Ot8Rs4mtn/uqNwuN776oudRlhqZhJxCiu0LvAsaUJs
9yEC5ba+r/S82XuXQ/chZZp6zhrIwNxPtUGLBJUqLorDJAWXmTi9RGDPMuZ8mIQa
Uq6pXnS8krljPlJaSJYmpD7i/6VuHRsyIg9B5oEetc99OxHzGW8wMX7LssTsboTE
DWkOKr+haua+SIELzXOl/YJ67szjF5sbY1BXdmYhQG4Aont1IcVVfeHgdFQ7Pfo+
pE+wBguqlKOnwYeReyr0qVxzyyBjfWJ/aIn+T6gZy2XStO1VHoNYlC88uDl+O6cE
/TRCRghr2zObolsoW4UUnOWY4e1QjmkcM808fg8pSl7enYiXJwqndCkYutAFuXGn
OoBpZQrePAr62MhyG2ONdOA78rYTo82a3C+jUBUo7D6HvU4KYFrMqCR5Ef3RAeVC
tB0DjdYnvmmHMfFMXU1U1O6F3LvpIzln88Urp3KDubn5V0cM+0dY7I2s0ZiTCLl2
B34PbJbI5BN23FWnFQtpkXI+p0Twl0dL7Q7YU4Cz3gynAHYxAXBZxUUQfPsFQQeX
xD4OeQfwq6sSbcDEVqSmaldro/jDMPG84O5yeanryZpKyr4Imk5wOEwZjvOWg2O4
izvsKgiMzOTtMbAzNYvH45GuuPkCEOzd5kN/15NPtxc6b4Hrise+7dk/AraYLTiV
EqtgbfvggbUSpzHFXicoWnBUgejHD1W6GJqzIwnmCidmv+csIFjHNoNxHT9o8qkQ
OokvWpLQuPcSIDE5ebwgv4tjPtqucJOFSfj9z98p/sU+S1FpSKbVonH9H0JstWHy
8P7OO9Ha572meNNHH56+6fvrdaftiyaTmQ92ePp82WNl4MWPCa3Akfx1iwGGdThw
UkPddJcA1NQxaKX9NeE3zWG3NZLE4UfoBbG2CcHm2Q+A5PmqR/HOZmgxV9HzMz0k
6TEOTYLg2WTSRvWos6surEvmq8FnN/tgdWIwQjcMvD0T0k7NYOPxKVZ4FYFyCoPY
Pg7n29LAcLm+2E9FrPdmuNLRE4s/UZdvyYpGAfTDwRhGXCVvPe5gkjgGLf+8Jz36
bKBZkgOwErsk57Wu9KqR2fYbXtkXEa5bV53nxuJQ7urGuJJbubbC8+u/C83nr+u/
h972S70MCAHsY2c+XyEuzVN6a7PsGuX5VEa2DJ+ymfst2c4eATH3PKy+QbqZ7FEC
FvvgIBdZFsVYoCn6IfbD8mjACUwJGpgjxSwv1P+RLLdbr9nULtAeUhA/MCRVuceC
GnFobWbkFAgYCRmbn/aOXBdKBBUkcibFAsA1KjWwOrNzFNQ1IJsO6kJAj58/tp8l
K9sXmRfMJ5D4dtKvvxW4VG7XheKoDhIGaNMzRCM1mMYCiIEdSQ+9pAfM8g0JagY9
FJHRLHGm9oLTA2HGmBTSyL/2o/l4AarDN9sLzJsHZ1lZutfX5D36vDdeedfeFwf7
pah3f4LAW+xDgC/tU1UpBAME3hpbfCaLzkeGhD6exRXB5WSmucPdtxTAqKsEzHAk
vzWO7uAPdzUmH+J2XCLB+9EnBaDFoXKiGSUB2t1v3Yo1GFHp5CEGF+/FMYORBrPR
ujdMxHeuXIh8rHAv9iuFgDqGyevDq5VY2/szFGy3gPgKqgYTGO0EjtDzrNXGTGzh
76dmAkCzWYEmIvnyG9pZhvVAc0mXWLdTie4oEUahI7BNBfbCLI+TzkDASRUlB5h2
0eoUhigelf8O0TJ7OeyNamK5FzGRGaJcuTSaKqXTZs0Ps/JKQCuK7e69f83ybL7P
mebQzYmgFKv3hMbRz5Rq9aI4Cz6CBcCdKa8gRbNG8FC2HZ5JuZfNBWnzAaovS9GS
51jWCyMGSJV6uYRifz4M7Z2yasAAnlP1acu+tdEqh8bcmcuKs5PmmrhNe4MxC1QP
qC5wCXXFQDWJqZ03dn5bF4DjXVj2y5gMkojSPo47IAjCaAXSSzjiWPlefEuwl07t
gJUPpiG9ZTumNdtEpjEooa0zw16VVHFFmfoLq81inXSEzX6PYTv5dsW0Axs5Ca0j
brAMMY3Q5fjWBw6GrSqlyL6FK8v3wMGVu11JbffSt9snmikTUjVCaBwvSb+skjaV
/zAvTc5m6iAHcS9R5fYO+ASUpZikbhfMtG2ROU/7BJqOGDdtIyQLcUlmD+bA/AUo
HmBHMWTutxza2pgoTys8ZEhNfVKcM3Iyfp9Pj4taIqnA26wDacZH3tFPLTp1UGz8
TCKyvXNNY0ndntWxdia9/K0IV3M8chBSunBLpc9CBue91c1B0icvo8nBPAcNH5UF
j7ICmbD2NmXSSc4MYuNHXsitAQsUAVe/xvQktjHLOz2Z2sIIEmGPneUkpRzWhwD9
oiwv/Nke3DZ8KnCf/GfrUmNGu+kDCzuD/lUhfquqBLRS2YF9qG4yQwI3Ta/o3+kY
uef98E1efHm8MBAgZSiS4HYVhfGJoR0i7Uc3z/oV/XgSCkoZbNeQee4l6t6nas/O
wUlfdFUv+N6eMxzYA+rUuG9ymWldHptBvi9zYJUtAd1rD3CY/r6tsAG3KsEVVLGJ
wi9hOZrzDplTxqA8kJ0d7UN0V4X4hIGjF5Gs8GuWp2olDFSNGRb8/I5lSZkYBAiQ
2sfb7xd3UkVXzD5J/pNtEm3/exJa30/PP3DfmEp/Y734YoQk5P1Dhtf0u+KuCFEl
DiIgiFxDDuXTTl6TJjcgHo0Y8HmVjnfM7HG9tw36ck8/jM+71lYt0H+1cqadunge
EcBNXg34lxozU2kvhYy52Co1SQFORciP/6NCgVIlgWbUidEk652ud2oi1n9G9T3A
GT6DCUBJdkcyewDyrPlyq1rdC2+A7cSpXHX58rSZr5MrEbynsLq27i846J3Lh8gE
J1RB5EHHFOSeWRdGDGbcALTt3iOyN1AxqvYlJkTZpb8mpx6uIf8tXVxVj5VelevX
nVUPWe9c9ydZuJtPZIXJiO2V+wG+C2fC5lHAhVxSXedFehGTxA0VBHeOZ6+PKoeV
p1LXDgeoPRAx4khiFDtQwpNKNPnEIbSQJgKAH1w521dBHz3mmdOvtt7AIwVWB74Z
RQAp4KLpLAVAyCbamP0mVojJvScuggbCu5yeXLqhxcG6bC/R8o4zAxlqaftQd3dj
byb4ZwvLF67hdQHeYsc5jXRf48WgPJTxH9No3qvWmmJQFc451M7vp2RJ9wd3z/Cb
8XXw4fm1N9loOyHmXQk4fJcA5Sw1Yau21x+OTPyVHYpT/IMjEp8WynbGDC87rxUd
VDYN8snsKPZklIMZ3Dekajhb1AHbWhMdSnicz6sHiXz3UazJK3PvXdelJH2cSCs5
TxGsZzjDzrk/O2o9ijgXFi4talvF++tBureI88oBdbLrmyRQjzVMGt+kSxR4bvOG
aQ0i2jbxnvB9jWmpSCRi4rb7I+F5fr8YSrYx6FStGv7zMHhg363fdcHttJFS4gTF
G7U9anxD0pkGsB94r6TJ8IDACtppRxK27zCPx9X77vMa5CCEiao2Om5Q0PNxgMKh
BUteljEYZarpqW9IlJviAkUREnu2bi4pT7sGKZtr7QKdqCAs6qhL3ovqHC3sZWNA
ImN1bg7VN/JeVUggnfTTK2YblQ5co1TpgK/JT9H8av5GPP/EAN/Vbw4yd/IR6ayk
XIj5ZZVCEbEC/vF6yPDFO1DWTEPBzr8PKwzX6iQ5VIJiV4Rbm7NmpdR1Ao9Tab5f
gxSEMcozuZyP8fQXfZSd4fDkOr614nT2wDiU55KT7EDEobHoLIhnlC/BdYBvZ41z
xCYB4nNkXrBdJ/G/Ihc5KxNDLNUSvRFKdjYfwsSUwU2ZhrwZT6iCXDcf6kqfztCc
wIxtuT0y2X809X7u7AMdudVtvH9d25ZqHaf+6RaFW1X50cbBfK4BQzQOAKzGP+1+
u0GQdqRkkhyawoJyK52G7NIJfrPeliB1onK1qsLskk0KvrQBeLJ4AohJ8f+Iz0bc
6t9RX4TlE4NMb8KP51qMauwckUhBbd03YDUXk8Kh7djjbQ45ArSPEIr2JDD7iGj9
i1ViShKLHtRb/f5VIDiVN0FXG0slzW/BwykB5ykaDuGEJ9SvPzu4C68AK5WvEvcC
lk+ZN5whSQ/mdGApFeAWHdLbLICKtcwqL/znwgsjLpJFy6zVjlwnyRD8zvhlNHgH
+QORoq3lHmfhV7Nk4s3RKb3ahLKrXGJnUBH9NBuXD3ruP4lrHQZyoe4htpENfCdn
9BsxOK6g6p5WgNNDCwIcQLRmEBF3r9GbgDyibZOAaqgZ7GD+8KBrLX+0vUSz+2/g
7Vdp6lj6FR37Vph3Yr1yr2D1ujbADIHCd3VAv8colQIsmkO1iQgBGJU8jdOFUNu4
tc8S2z/ks1gdPpY5C7c9OjViL6RKywFIvuh4Jl9UKjbWhTYUUHD2+ZBCzLiPcTS7
ILKmErGnnZSns/jctyGtNYjjaCcofk3yNGE6tdbdGEw9Hw/qnFlTjn1Ve9+quFz4
UTkWs61820k4xzURxcd9KXzxF4YSqjdAq8p7Z8lHIU3RoH4UnuaQQkEs07gVBJr3
TVZgTGpvFZWaZdqktIecmXUcY6nriHGY/PSARnoj27bXDw64x8PYlToPYTuJwmWN
IgFBZEKMspIlP6d5aGCzY19wVify9RHDgrhdMbH2iFb6uLQZYrC+iDJWU1qHZgvB
3S0Emi0l/jJyxUh20rt3X4/A0X0XyrHsV+KHmxnK6qgZAfQeY0g+yCzLHBHJWm3U
a84njAYuHcL8gtYypgAGImtGvFsk7pX2R8XRXwykAjTOiCBl9ozt15nQ/z8+98xr
hfVj0UwswTBgyMd5liKHAElN0YmYBF6Xrd++ZNUCigL6D/+x7hPKwVfSmMKsSI7W
dMk/syFTVEJb6t6dWf0kVD2duOezoHCK6OQ0aSjrWdJzdl7RiN3bbzhWTKWXsYds
pFoVKmB+sstRdflFV2s7RMBdpQqRypb9RxWE33G4QyGgOsOnZsEixZk4uk2ji+ec
YVhSTxetwfBFMYfbFpx0QKr/nRtfS6fxd7iko21pqzN/fvMrcpOTNEO5hJHVXpWH
9oScnMBcKmfiOQnSLPlTA5cpjqAwlK/sv31hAY1VmrJIZ01OVnetUO3CzNPSyK1R
dWanGWoEroUcQ0pQlumHOuEn3hfqZvXNKsBrQyN4eqYzTOUBzXRvX4djCdEzQftJ
x4xZ07wDsu9uoc21Blo8L//YQhmfO4PDJE4K0NEJFI84Lv/DIb3J/320eGpfIz74
LHtO7i0LL9vpx+mUx0XXInoZk7h3n/JfoXLkMGIjzr1G/tNb3hXMCZdtsmolUl14
y7vkZ6ZCOm6FswQ3y5D9JWqTiSr8eiEKOEMx4NjxZhVXZyELwcjsR92mAI0I45wK
EiTq19K74ivq9i1has0R7pmM7IZ8drdTEl+DbcKCPYi/JZ2yhUKuEEPMdNw8+5yO
JAxh9Ug9VEcnwkxoN00bbWsEuAXDQVOEE+16BFPbTp9GtKSnWi1iXhBwNGRA+5EH
mZNXKGCl+2QqVRIHEscyuILXmW9KiOVIbHflTE8/1f9KYdzfNuu/Tbg+cYPkthyn
c2hfgwux4aZ5RXz47VvU7YN7FJNBlSnxMc7aVsz+kQ5xw83bARY3RXPC6xyGE/Kd
dFQsQBnjREQYuBdq4Ew92l1OrB5GKeCa5KAJn4EOs9ZYGhHePM7D8IFJEgSRpCAY
Uip+EbDJlfExgE2kavECUE0TdWwPETIuWmnANlKHpCLX0HhBxYft7pKR3Y0CVvfN
9r2z8gC82Gnp1mpXac8JBJqMNseZl/mRb3Gdz+qMUYU7bQQtoV2U4ax5ke8nJBTt
19LCQAlPD1hixaswq+hLkoV8Ywv8PsdpZZ1WitYhZkya0C7fmY4wPQ4trtYToUuy
noWTrY+qtUKdjOqGYuzZiBAi1nIcnEs6daMP1JGSF8SVu/WTO5qvI/z1+AZY4FNr
979RJNgNvAA2pFXVSaayCc/JI0KGcmb5l9W2WvwTQlHsZCKL+rRhZo+y6bz31vDQ
LsHwsci8Dc2y24PxkbIrJ5QqgfA8rR+uvcFA+6s/MUF9d0mxeU0Sgzqs4Md83ZQ8
4RaPA0EnO3BZH2mjo/6YYK0VMMEg9PUj8+u/2cmyeVQ9U2nUDyTlxcO+OfazsWD/
lQyCd4WU95b1BMFby3z6vlEM3fEe1hDpveQYNfO73HLitvh99Xzu2MQJQfBIME8f
6Ut/TciTvLNLwod1pmxz/l6rUl/ksawu998N5kk8guYrDPd1HxM8PlhGu74BS2Kc
xcdAawpBezsVvtHaQF8clhR1eddER/Ruy8K+Xci+0LuxpoY2wb/zo/M3KyjzZ1Sx
ywU2/1H7LsEcgzmRPKihvj3RhDzcQ1rG97ZaCxsAr0WOqkaEXmQO+Y4ckAj0R++w
zYFaNu14UaCGpKxicHqg+/Bs8DNqNFwxQ+NA8nlVrW7w+wTNQSkDupY6GPkATw8O
KhxgLdVIZjepv4BYRh8FGzJmV7vCCGPgKqFP5DSyTZ+XESST9TICrJDqa9y/TgiK
iay+XgPiTERAMTFgmiK1IotGuYD58MVRD394sdRgeQ/HJwPFs2JWKVBXmP/gv5PS
CZfy63tQv3QVDU/HVfJf9++nO3BTGVUyyRieISt4ChurB7cBnp7MjcHmq6So6QPu
Oc1eCWjFkFq4YaZL18DEVioxzqaj7DT+C9nWJPj4Z4uFnZhtJqOOH9d4v3Z2zp//
6zs5+I3IIHWohg0eLpJ6lQGVn4qVLlSZCjfIVYOXDmir1lZmqXzvLQQWJl6hGd+w
828jgy/opeSP+dyo0QsGp8a7YZWMZaeI3degj5Z2NHmyILu3MZRkRCb+5mSKSwFL
7jo4iLns6tyLvRpTx6R6Xh/WLkuXB/iKWSA/suUGzjgf3DUh8uZTDEQ392/3+aRy
ZExB6Mt6fcDYAZ0KbFMmNz0RmhciAdK5eZ0eM5imXpAZde2knsPLiWxEe6lzDTPG
u28SZj9DSiahTt5Sd4/VYFdbI3cZUlq7DysWzxvkoW+2gSlkpUyQ7pHC24qyYr85
B1qBLjkFrbbcYMHXSTjjeVqssfAswMs/+s9QjMOr+ZHSjN8pq7WIMQ8qNE9Q8Eki
fQeb+dfDNTzKeI+RGhvGVh5wvCVx4N/uLe9WF3lEbkrnxk/YRJtppgadgMPC0O+4
e0R6UIsOt/Frv2nfENc5zSeRXz1a+PvOxthPwoEfPGB5Z7zdXlLiE19g7W9Oygpd
UAHFADX6UDwVci/81gp41XfU/Gbwdlbg+gfgUzEtjGJ8TMha3mxUVjU21sYHHm8/
gwVfeKtX83Z4J4QAYWqlYmuu1wHGrWQWVDtky0Vkdlcz8iBOllzFBDHBtxccp/Hv
7dEUJqRg47aPMnXHhO4YgMZ28bO1OcaoHdWc9pMThrSzXkLyE4aZZYo03tcKgBDr
1sP12UfFcLxQGjBCSDC19eOoOPDGfCrv/D+TNg2VoZfORfYEg/rfvGFQRtLvhHeR
3vGTgJqNuyjW+q6IEi+u95kvbL7m6BVxKvdpYtDzejef6A7PHg3dva7iLUDLDplq
6Ir6qkv+OVTgRztjF2+5zWH0ZJnZ1W6pLFWcxz7cgxDIAMdYQLESN+deRLGB9yRu
Fngv7yVduJWiVR6gvtuvSfmOFs/4H95TnjhADAwF3wbxaUN7JjBHWyE+sxpQvKYK
7ZpFTwNDVCOKC8I9JoOpWqYzrXQ9mfMg/7255toRzqwYDgxdjW+DqQfaMxusHa46
XD8/QUeQ4MUyx6vi8c36kLYFau7jWeESVBCeTCa1y0Em4SQzArGRq7XO+7R5KNCW
n+ah8YHXXoyaTNXuwNWZLVJLqj/hUyLZxhSzRAd9oUHFLj2v/llgCCbGjtz8/Gfd
jfMYU3eaFA+FVIlf0DqEEwpqLgGxXMK+lyzCTh0SIpJl0XbfKBCc1/5Y8EAAMBsM
ZhfU4uEnpvtWNXh6cWeyQQ2FuZf4yg4Yg8y3xZcFZ26mFDn+ZB5yx1ZnPQWMRw8W
dW9SmHWZAOSxijoCvIwTULwQgKqhuY4rd1eds8tGQ50OJDWQLFGfdtwmx6w5mngb
4U/O+UerUYs5SqS3D8mwuZFkXGpe2kwakmRBU0uca6KQAvbTNiyzoszDQpLmYDIh
2lEFu4IHQ3F/QTLiRv49+IvySamzZ/wN8eYlfnuUFpdO6NEeT4Y9Qgo1PUYt6E78
8YPTLhJYvmIBCOStQz7ni9/Qeq2up+bvvMnGbyMUPpKSmN+uvHnATnPTZXAaXI4C
R3gW51uUpplw97DbO9QN2TQvLSTf1YDM+Rn7K14+5sxVJVtWjNim6+mPSDquZwpO
+NYG1nF+Il2uLAyb41KVaWwpKxUmvoSjyRtYNIWpmvnVa94FaLKD8l4XtOzqiAiN
LnMpjqyMZAa/GUS5irii0kTvZvjiqXIcptap+ReIH9AAYEtgVqLdDDe7C2Rg7kWF
57/6qe0CrMcg3braRNZUtohIzF8ecdS5t7MgFKCyPvjH/x3+NN2E49Sh9aE2KOht
w7czAhLQTm4IWLCqwzLmvwscR2te+RDnU7vX3vWgAT1v11BtqfpYI9A+YWBLs55h
7Rk7Nmp92nLJaScPS9PQvniDBv1a+4ZUnrRDa9BBQgT7d1idl/uMa521hYzU5qX5
ZjhRWEoIKR8cQjezaJiko3tI+Ih+bKu3qoqDgN4+45pCEglFiN2aUxeadSD+8qTu
R0MUhB2MBp8RmW5K7vilavhv2bCzMsC9T1o9bAs52BZ7XoaObpeUXn01CTNvXLRG
U8z1vTRlmUf7N1X0vOaQjpX7fnowd0BuLeAiWgiDxyyz92qZNO2PCVdvz4qbwLux
TLwKSr2IXNXTRJv0qtV1rg56vo9X3lLimOvHhivU/+8pEXcZ5EUDmjG6skaQjIVZ
t2Y7k6zyOC2/k4dZijV8DQYYkGvSLzX0eMOelHtyN+tT5i7SdHQjrVX+nRhmed/M
7Qd4LdbPUyPmsI5WeI9LeccfCMTa26G8LcyXIyDmMvg7uJS0CSj0DCKjXzSeVGt4
ObD8QmSB1IQLVrlCZiDXubmHgHBtp26IbtBU2CsZLB7X5hLYO4PId0BgTuWB4sfd
29WCOzGOn/I3HjH+YjuJm+n96bJw/L1fNpGi7xD0oFnoUTbAnci9M428H+eyrApw
Z0CT/gEhWOkK5mkaaXa0mdMtDPwxYfc3D6gyjThxQeJVAE3B8HHxUSvp3XY2J89+
yCtrpRwwfz1WGRKV/zHdQfLjI72r39O82hPb9C3OdQCjqZ1IThmpXRo+lWTz3GtS
coRg4PljzwLpxto8bBKWNoTBhe8FfvQ1iQQ59pxnQxiN5oQa0atnDgo9o1NxpOQK
EXvIsfpAoGy/aR05y6eDdNAWhnoYNQqrzziDyOoB+yeyZn8PvV8DK7iTFpM14vAu
Vp++nbu2ku+87wRs52JouTgHy9HOkMyspKF2ZaAkH0X9e4PG+7LGWER07DyX7307
XP0+wpBiGQH4gMZevXN0JccaR2szhfUrsMTyNARkCr3AaHMBsCiiQnh/1VP1dvWM
3D+cVb941NYOqEjD7DwQWjH1TqjbZGuqeQwPuNq825h2SupsioHVAJedP3ZlpRz/
d8iZerWXrqXxUpKbGypQY/z273bzM+mgKJzdh+Xy+fBj98leEBrG1eLcDH/q+Bn0
wFmXx5NHxr/yY5kBm+Ai0/3ldOf4vQfDvybLDKcA7qDzJKHLIsEnizU/eETOOf6b
hp7dVyYQkaJoLQchvk0phMwCvsZAeil/Yk5v2m4yk8P5DMOTGpqHlatgcOgDeqPg
HW8x6jEoJlcSZOKdg4o8/8+X7niKPMRF/UhLaJvsUgpE7qQUAG0/bqD73FE0A8Dk
94DELAhjrRe+J4LX7Qaj5Dw0xvTLPjDZlVXSDJLglQ4jo3i4/wKzP1v4LTtvBSWj
pBFTtc+00aOoxeAlp1gDEsUNCbLzM6QnDjg/Hbz3edpRefez6NW147XL/JB5Z264
YNYl8kad3u5XS48qDWFhjvo89VqRB4MfZcuKvmAXnsiTzXZEK/kxgguwoEJiiik0
r64vPhDo2MBFcTPuvDsko+sjc8HXWuhcYSMGUG4zTTzEqeMW397vn/HXQIXCag+O
ero3DARj8xuBDqrFj846zjJTroVvKwws01wVPSVcxdxnTeNWfd6fpcQedeJN1ec9
Cs4kWMnEEsfRc3ZtAyMJ//L4r30bCrzpDxYvcOnoLEfSs672sgcGiEarYnQgyEOn
f8LbBmeOp8HC90u9FHfAQXmwg2ORYQI4j9xrUulrNSr+R8vDPwTb5Owwyt9lR9vU
ZVzXGKExqtAiHPLx9m+JBLm+5EhUrZIXIrH+pHvjZDXb2UumHrZraw7u0LF9jh0j
igEwrvXxSPbywvCtcECQom8Msss0Qbgoho0VPHb/7ZaVQ8htQW7z5aYpdtW8tkB7
xdqNUQZVwYxHZJ4YfOV8vZeIacE+c+JUAOQn0XCkL+eBUaXipYOtOALKVrxHWPtf
acrVOFbLEXdAzZItOt86fAv3Kv/pZi+j9MXXTjZwYg1WE88ZsEWbPl4BRNth3hKc
xL4qPtIGrESQ9x7EuBnd99ZYdvGYF3sM2iVm4Mp6twXChlXjUBnf3XCoSsg8WXn7
1FI/ohbtNM23rqwSumOTluFmk1LO4F5oOZeFkG3gHDnqcfT3KqIY/mQXPNWUtXAZ
Q+Fklh0KhCP3zl/FENtt99LCN9WOeKTAP8r5QQ+ZSy88OGD2WwR/Cz3IsPO6+0aA
3qQGx/77kbSdz7OvI0iBuFYIMdz4Thwo2JiYx5Osd3WuxujLiaO0igWys/BpVcni
9KGVhbHEr3ghNuyPrJFP9kQyn/ODe9eA0jzWsMwXBT7aZcpTfryNM60+bTmYUYZJ
wq8Mo8i3d4hlNM4rlpsaICNus7pa5SUa9e8N0CWMaYKTCbC6OB7Mb/ibLNYTLxbV
SR80aSVdJJ5hPQ3mrUkS7Fkb2mtcwp5UCi2BOFEiTfzbsRYGPIClV09SeYMPrMuF
CKMQh8tFi3vYPBaPu//0y9OQFZp9RP31GOa0f6ejkaGeKzt8s29MjHo4XhkIwrbD
1ktjG9+km13pDqWPJdO+FIblCihDvrfSA4+PpwjBeMiWu6ydD6OnqVyhDWe6wY2g
c3jInpH5KHVklLKSKZZKVhxwSm6m1whgqSGhCw/JXy9r7OZF5FGUs0HP7hxYOY4S
sDBl1jsK56M9UqDzA2jBkyfoD8w5AvCEWel96aKM5PUtDs9D4WbZyxfmpDkJdtUh
wHzZE8hJJBU5EY0S70svwo50T5uBmtodE0MxzyOKerTsuod2SrxGMGpc5C+doaaR
zOuL/FNAhibHXe9vSl8Qu3Lhqr0uPSFs+cT+BI+1b91KNPbI1KFjgozf9wL8HApr
pCoL3MnCpdr9m1DE4dceuTzvza00hioqv7UqlN08wz8Xx7Wt3CjkLyMGKA74vo2Z
9YhwVgXxbcunO8E8pHSo/8zKJCVCkghSBsarxXlmnBBuMwHSl2jtdwoFqg3gTVXp
uUB5bVWsTddLN8NvGeobUoQi+55NNoOujoMUJBgUlQRN753uXwthVOMBr1ZtY/HL
B5/EKn2EoPqSpTywfpkP4fDErRt8lKPm+M55lYTcva17BvUOQA/JmxN5ySxg1fco
yzS7/KxoF87VLFlD5Ah9XQ+iR0M4gvCA0vTdX3JHgeB8bIbnI9UztMl2dW6RVKfv
St/XsJIhQXyP3o2xAu6dnQiJWIB4wnGwqoH1Kot+Hm6c4dxJZtCzONYh4MJA6pUJ
wNVfMHuUnzvJwqF6RaKx/IKOsViv12TMVyPr1jtHY7DtJ4DeNVp3IbW4wWZqsUlA
YnAHNAdQchLF0XsvbQ2xfijK+h2HqoOvFL+yhu83KWI1W+L8XA24gXZGYFzRC4dX
iPXWzWV0tfgpiKSac+t6Bu/zHvMy6bRQWKbCnm60io8mIPObYPikDpyk4/LA4ACo
VbWwll2bOU679uAZoIdQNkDTUzrOvUeAubzmH3OJd5D2z2+F5dKIKvAbQ/iyzMhR
oMhz137VYxU0MEGLAnS3D3B5nGNNr5M954nwBZ3DtKUBFI7S5a17wgqjRNmQU3mS
57LVk551D4s7m6p3zZBOV6TkMG+Y9nDdYTXwNOVi8279xzzr7rVZgW1KLrWUbKck
lAnpF2SvbYa2HKXgQVLnt+wOosN+ZfrIw9dDTSU4ozRMNkZS4jlC6i0utcKEBcxN
vxRcb8qeCIaoXg9kKmg6syVZiqMxf+Jw7exCneZeSsMSMhdmbstusgsXcKzELKYB
JfVjVmv8i7uMZkWKLzYPKLNph21/GY4RvQhY1NK/vPiMPdxx8z+7pBdqdYHT0Kie
HcvUDBXf2gFB6DKthSv8LcYUOoMfGkPtxNu8XHWTTefaUVQCrxg+8TWDYN6/M/fo
+KdJ7hBD7MlRsmZeoihTGOJj7+hWgnSb8KPyTxImcpciOCaBh+q4VypcqXFV8aCl
1NzbD3rKnUll3zQefKUrhlvzmP6m6L4H/mFy732afWKcfl6Glb0tQwqTtVOITqtN
GXVHFxgwtx9iV27EU8jfi7wjAkGC5K7SEncJRX1WFwOlX5xp39JktOmXoSJaEpx4
UMXK9LpElDWqIwCjRBdct+Uo8lUrqxZuzmWkTLpTkWkKSw5j+ZKfy8SToVIS4v9i
AG0Kk1pZ5A3ABo/KtHrVz9VTl0yAogsQyU8Zz+2G8pVUmYEYO02TpbCecnsgypdB
uKnuFVfCI11wampCaSkJro9f6ynpe2OmxfPLCddFOgmoH6V4aZOLw8Lz3hQLEOgr
4fSRrKPyuCxPvQKvxeKotlzwzZjO2MsTvTh6YFILqP5efO+XHN8Semrdt3IyBnZ7
SrzgUA/bXXGh5JmOSOYExbKcGhEvFuL/4phunoO6iSDaFinraySdz8pf4a+VQb/c
Jy0CWG2Cosf+UFkhpkPe7re4uVWEs1V9ExnwDDKMxjA1nmGHHvDm5n8B+lNS5Jnm
bYI7LK3ItuJR0JWuQKbbYWKyTQhYHkqnDISgwQCj/mluKiiPW3y882W0KvxDF+Qm
TXS0BdYoO29BLJnCpbGSMItDKp7/zsG6eWPeD+2LJBcn2dMmw0kVeot4Ghx2Jdiy
nP602LUywMf2UHo93ttH1Kf32yetw5Tk0wNPno+5k4jvDzMW8YokY3JntfQif25o
PyQ6PqQHT6YPkzuik+HroH0QZZGnlhGYz0z3B7p+6bhebOk3ynK6MZH7F6q27gP7
yhOq51Y/VyHwehNC7ior4CWIFLLKcjOkxXsFw9cv0u0hRY+ZZzu2Owd/nEr/HZi2
8B7ScG82mDGUYOGFbOzqC68sBaX5skyDO2WIHMMcIGEHzvLkI7ioj3fGQ/FnLK9V
0ARctOPEPjiDsaUXAaa2OAwrgJAIQ+4Qp8Bc7VKtBOSc0jt5k/HfXfhjKotz1nXZ
UKRbq9ZIT1SOVUcg6SypN4uHaaoVSqLljMOSpBIDC4a/U+T/BDSSdt+vv1ivDyg/
GwbpKLKaSTQ1uHKkoAZlY3WeUGAcqoG4o0XbU0bn7ZfsolwxQx9O08xN/8ncekSh
kNBY1kaMlrWli2criEvLizk0kedcAaREwd5KAuj8XPFqrB/Y9VPnlAJBRGngYhpA
dDTsyLrd48ava32fQzp7ztEA6yBzz+snlE4y8GnUWfNyFoyfeB9tXiASlov+keWR
2uhln9NQLg8TjJH9+ucZ9H/Zz7vZaoDBcJHN3YLKX8z5ARO+miDcCgpp0cq3CqvS
bI28tCOXXFNnBXU8nrsGMmYCM9bKxIVY3D3bFj0DwVxCHUZOc2rQYbbEhHPKf/Xt
yvrp4NjwOpHj35+DSzm3zY3N+QqBvD7NbHUsQw4inc3z+i7t2jYeNJAhN0OgoItF
r28jmfFJygXl9t64P+KmjOLJZybMzJzAwokBKUrGi5HK3C8TaUm8j8hulsSW3apb
zda7hokHAr7JjmumXBEiQTIPW7PqsjghScv/cx+IFtGtKRQXBYXj3UA/RPpQ23CU
H7Y7KDmc5KZW6/odjHK8Z9ZU81pOu5Hz8EGdwJxbOd4ztR3vI0D6/Ppjq44uoEIR
ooNFvkHWbgAyREEg9PlAMsqyj4Syn64zTkZH65etUdtoagmrJxA/WsjxrQXnDWE1
nbx9tQTSpJqPejgB10eH5NDPmFJx4Di39Shfis8fADSwHRkAW6bGQ7UGB/S3r/+S
khqFdZ/KmgTtiCssRHT7/d2BYVpIUFt9ts3R0uc/FqDGiCKqiFxR11INmtSQQkJm
guYOgk8WJy/eeCrUPt5bhMtm4CQCDuJYfzv8jR9T63qdYQan2LnX/RQYl0zg8iL8
4g56UAXbjrJoWw9kemFLGwo4ljD92iXfFDFgD4nWO9lrm6fYI3mBJhf2Rlzp6+aU
9Jiia+a/wSKF/sawEs2vakwY0rSgs1q+F/gs3i4SAI/wF+VbW7kHTCToJVOqlQXh
24tX1GBMDOcAWeR4msLvXahMAjvrxSC5z3n+tAdASexOTZPLO4E60YBkay9eTUVI
w+xfE/6qwxMT71oV025EXT1bUtbTpqhrAud0XwE65K8CUViG7CMX0RtUDRpsZ7mh
zsSrhWj7+oP0SBV1ozCaY7AON/fB+I114MhJVBvIlmERhDXr3vI7lQk4cSjxOy09
GBvKsOs9Aqfi6KWtalrY/EpinkHd2HM6Ks8+oc6YsdXbE2z0Ed/EeQp3l190o9wT
+A0Ojjam6YYIFgoIEWSGJWJlVM1at0L9IARQLXsLN7rT3JLNscHUr2Zgir9iiNdt
pyZPXmff9yOEeghfeTLOGql+XZ+TYykrkRHwWdjS+V0HrMz+6jK7WQXn4xtAcB1g
2D+XvGRVwulhNdlMIEADtIP/ZBgP5KPjwabim8jW32FhszAICnr8xjYHvjumosgO
ahxOKNYLV3HdvV5CLMZ4yvvrC18XV0/Se0xZr/V0vpIJVoRjCNF2XmGdAR9YYhnt
4lnh1Fh0mt4bVdH1N5/WfBYv9GUzis+1t8nsiFJxpr2J9sdkCQNTNwQk7nMoHKMa
CG2qKOFGLCSCbwrWUO9vIH8kUeDWyqrBQ4djfzyANv8yvGOdS1gmaghLt12Q8dfz
Yz03kEzLsNHb8x+LHh/WAqbgTP4JsMVt8TZrzHvwq1vYNA8DtzMD3fnfmbQH62hO
snshkBqQccVS8+8QtpveVSS9aj5OrDhtUuCDxcT6R1Fk3pxx0oBTCqEO7566qwsx
IgkcAxWQ4C/iCgaScoB3tbvH2Be0gXEPkkAMRNAR5ZW9bOEBc2qlHHgsRJP4Fxvh
Q/pOVbv3gfNmP3eORF1+Gr+TU0idXAzk/f1+zuwVHuyoIBhxL+OWMr1fcoEkdDPk
4fGBudqWSkmds5X/a3D1TNLbpkGeIPMJxw1suQb0Vp2IMQrRmZogcgSUXC7J13mV
bf3R38sMPHImwDH0z9PWMcLyevMS/ERP4PXC28x81G7rlFg4RBwJ56yifEtz+78N
kO/W2V3UpTiLBeEMv33caMm3Ec16PGInpZlhoX4Cwf2doMAk0KLHCacPM5OrFo7a
PMeY28Ebc+i5Cr+DP6o9epz2D7a/ALbyPZhLF3IY1MzQ59ImBiEK6NW6eMTYMDdG
wwe47Emib6G/iQYDxREjv2hdIkSYM1eqhYxLVZ46Idx9u3QA9KABFwXpkXGQTK3q
yxTDUHZLQY+eLa/LWfIFY5CZMZp+L1CPIzLgnx/gZz2cfgH46NEGgEPqtVjxy47P
XL0rHapmmprwgtcnSoHnkjAK4aPnVN0krKe+zQMcSF6wGl/dWdpBhmKXs4IT4wOY
8cvy5OQ+Wg1SKioYHb6pcD78n4dfRTXmGVPi0n4FwgLHcgklFmBvy7RbteKv8IG/
6pItInHSLHiH2d0FZ3OAPvQRUZjWxfTTo/ZQ8bO/7G4Dn1q0X6swt/B32E7nCvBs
TFA+AVZuTz+YboqrXzikRgQ/H2w4FaX0MizBnLAxwaQt20yCV/qJfGpEFOqC3jff
KIN6yLIpHwGnrBMRr1TTmNOCs/dO3TspmM0nGKTSKz6Mpfh3IEv8J5FBbcOPXwpy
1C5rQWhRlZsZeQ75P5F+rLp3tbd8RMA9FzJqg1MfXKwYz67UKycqrMAw0Nx48ySz
kFvchshyuD7oIQa3qFaFDDYdvQxCg+WP4+9EwEPDrt1ukbn/XlO0WQRmM3PwkMUj
7KTOwND0ypcdTdRn/JMG3Eph1VTenKJUGP0LQBqL8f/xJUQz/3ZxIpw0FHRymVAd
Z4KdnzGgiXQznE/771/ylv1sbkGwS36OikrVgWNBakVlmCBCumb8XzC5Vc4AJFex
/e8tPzcLTGwLWequ+jZPYj11ciVZAA0Ro8UyqoU+Qevb5qU2d7ta2vprkYawCUV3
o8KJwMP1qWriUBvw2FbKd9oBWarL3WfCJuDAQ1uofQWWyD7O+4C1KNRLXjEZD4NJ
LdPUfr+UIjSnDoQyPW2MbodghVo99J+lcVZzE3JwmNBNlZdawzc/kDHAEw/ORwtW
gq61d+OUV8HfzG24ZQ6ZDSOU/pvdL869+HpSVkHxZZWxEed4M9/v5EhQrdNsybsY
ovFp1Ih+4kuXVsmDrr3m3PklcZSWtmIJ+4zkOX/1FJgiHAIs1v9CEiUh5ODLtaKL
EXBQAUa1pFfILIm+L4tm+6KRQ64QoiE07mL4+AdaAwCnhQ8HSz8qGEQ1/xQKq+jP
pu1wMEC3HWWJ5oaNiMTHAn7JFGAvlCaO/Hz/yMCqpHJycK06cloPHgaWe4vhD0pB
XpDEyZQ6b3e2PR1QI6FFkdTeuutv30rpW3BIqy+a8BW8nwzvr9OUZXIFvXOfzpU1
9IKFvkldIZGnXe820YZVikz6adM4+jvwEhUtehXqIPwRq+wIIerLsih3XTiwOJHQ
mXfy1zpFLAZOuuu8Ao7aGnR+Kb6HBcbRL7pQuXPqLIJ8YHWUNOb/8p9Wj3qTTQ0/
y+TvRLRVq6LTztTt6Hm5lMEpT+ZoodeymI65y3rP0EVoCnx4K99pm3P7awlwiNrx
oJ3GIKBaOLdy3Th0FP23iqYOgvuDjVqZoevxurh10wanXDu3IFc4NopP7uDkK6XD
SySh9C3J/9keTXEDTiMMNEVAo2OxlF9H4v9FLGjsY+k5Q/7omWTkRe2ckTfqWuGk
l16T8m6XQXbrMQzEY+kw4qaxXM8tZzDQ6cNflgDPEu7poL9pTkIHULp0kifqpE4/
Wbownu3w8jZxOrn6JoW5AHtbPBK0Rkpt2CXnFB8OxJlvzSrrvL0+W1zPPHfMOd0b
HvtKbt91BhJEHIPxWEiVRnbOqCS/tsMn7G0rH1QESQM4EOQePxIklCIIGYWqB1Nr
Fp5e84UQlMbwa6dc0IKNdeacIyqxRpdZ1AZ0Njs9Pf2i2zMxa3Ke9czBweoGEPyF
PelNQ5M/h97ufw36Z5Ot1lJrWD8Nt4o3wSJOGGy4+f53rXc0rNSAvydltb1Uw6cV
wSB2ZmFsZrS86gpnT3lFpBavs78EMWsvRPbQiZdFBeuT7A2qjDOlr7cEYzZ9YMAN
pzTJWeT+Q8p0GYfpTgFebrV8A70ldzPOvS5EdUbDHGocnFOorvSVOqEezvWHQLPt
iDgjJ+KmRxU6Vbw4HP7nt9f0XDNgQWTYYiOrqf9bHVaNt971/ng9fieVFwnZJ23p
oUnSL1sr/YM6adfeOMD7s9kK68qTBQavfek29P7+b6N6LzRInayeG2i2M/qOdH2F
gNCIUE1b2B2j+ISI4cvOmqlWwsTO8GFq5KhtbxiaYlP8my/cqhT55i3tbSPoAzyH
LZTfoEG685Dy6NGY2AZF89jaQTeXPQ2F6+41zFqVALrKimGjE24wPvUthS9/fksD
5yEEgUgsbW0Re7yb/F3EwEk+vPcafOyXjmYxLigVUGfSuuoBEZk5rLr7/dt/kKhV
Stz+ScD2XHYPa8Mf42ucBBluE8NSZ9ha90eZNEe6ArOz1WO/myAtAUjYZAqD1atP
XGrs3/jQBIdPUn4Pbv3dLeFSGFLgMb0xxhr/EvYloeAy3NCSPCbRokNx0LDqJhwZ
gjI7/+KSbbT7pnpgpLfdPzpPHSU/vjn+g2/5WaC2oNXxlFVvY/6xwVIiVf5JRYZG
grn9zoEH/AA+8muGFEqraiQp4ZZPVwWV1ZAlq928DEgnDPmWbipIr1Ea9w+AYdLW
37uA/YAIlfIxedtAvmWyFwQFxpM1KV0on4iPGLeEH2DhDHt6sOUy6aEf7B4HjAcs
NXL4IcsYurowEPZhNA9XbiwB+cIz589Yvtx/bwZcXBjn7eJUZwJN1UqDG8gcn0Xt
4Vj/fbmHPPWRHr9g/x6ohUR3SyvReHRE1/nmVIJ4jiCxXjh7jYq5sMydSZ4cPJUb
nCUw5xRi+XQ1MPhPrSJL/zGDXk0VqMMts63jJSRdN94SKhLuKBlkeXjz6HOv85l7
QEryUBbCrvANfg84C+bqLzhrK9uTUhEXH08kQVSVXJ9oDzfn4Rd5uqo39SvNKGp3
f3yfxGw0xYWkmSxwhzwb9sFNgfV19QFo2K0SvF98cxqjUHrAKV/Ex+nWvqZHwg47
27z+VR0wfFpqvzlkaZGotCdCQ0nj8tB8rJ2z9bQ1zLx4vJ5K3TsjSbxlMDUsp7D8
QfUC450PVS7x+u5j8es/DfcN+lFKrK+ACZQWXqJoGJz/B3eMoSkM1s4bLCslD8c6
EzB7+VQSExOyUFEYyd5ez59QkmtgUTlIXIWXtIhhiI9U0ZjkcK5d5RBAdXTyVVR1
3ALOpFGncUr697bRu1tZUum+zM3f2PYJctgJ6bgw1u25Skkjpz42Y9wTkKCyK9lT
OYVeym+EAoqHGC3rKZpS+3JkxjPXR251iXMBPGs0SzUBLPVQKQGEXB1XY2lPVBHu
5iUIjO6yXuJQGQzmD2PeEOaWHLWPraYLnATu9jTz/qVEBbOx0+A9LloCXMDjm2df
v4wTwkyV0jQEsWlUnpU+dzF9fk3IJAqXw8m+ae6fJ9mF6TRIM0+ZOVPAIvc+M0R1
/uBtZ+9uznIz4Dh0NIL2kJpNoypXho444S+/e56jKXDIlc62TmQCGI7bkmikWeCa
Ujsocruzls4KKndQ8QPNktF4sxDC96IKzgyHi9C9NvtNkxj1caMFv7tfUewlKa8w
AG84Ow0iWK+JaJ3S9YoFY1GYRwUt7PGL891kiadsDYa+ku+OlInNumesBA0zj1eX
rHPjym7KkZCKkO8Vm7MxY+cAVbix0tsMdp+g8rhzJlcjwAkwYycMK6CEm5waMYWn
/zPmJ6+P7gVb0nIFEDQb3FImSBoSiqEekudOZ1A6JFSqh9bNC3W9yOh6dRlYcbud
YQQaLuTh40LfGGvB+OfPDBBaUX7K6A5NDAA6zL2gMxJN4fcOPDvjLMPdwYwT/4+n
AvnQ+g2w3novWNJbITWjkPd9IPXdnercd5/oUcV0+I7GhcZmcHB+doFpgzgFr9TM
JY5Fz8IfoVRjCxADYMgOjkZImRHgQXW4JR2mKW51+JvuROEU/5hxRhVBb7qd2Z6L
iO6oASXlPyWsguSYPUgn7wk0SUthIucrRMNJ8PPwxct/OmcpGhE03ooKK7PiZFAk
eelZ8+hReniyNE8aP/pySpFYvufHU8V4ygUvelvzvDYNguXLPOi14PXPYkO3quYk
Gdo7iz/pPAu87wKrvIjAFqBstrX7CXduwKeh44lt9dhgAJrmX3XArReuexTLK/jC
gTA/EgKGmzIEkAwfc7ItSi5tx+n2k9MHK2cqMwSYOVuGJuuhvWlmgjnx/LVr7GTH
RCe5QTQN01rr/aNgrWONlYo9zRMBIS9mJWFBLBpaRxWsidMJ05gPAOKivSLi64oK
YFxnbhoZ1C4MrJTnmksClQ4ljtU0OEQjraMP508IEIe/RktilnNJQf7rws1u0iXN
3mPdQfdc0jvMn0g7+x3aKur4SdOu/mPU0mHfQMSTglAfupdu6lPxiM5YfHFl261X
EH4H1sNNpQhJjg9ozNSBb4ISZ7q85XP3eV9P7oCeYyqshYUH6wP3v6TqDzQqW8V0
SThjU23tkBK2ItBK74noL4GDuiM8Zyt8B7deJU3SdBzfKt9sBa8O6vVPWVGsI0oo
VmJMTqRvGiZ7BiXwwQyDPl55yzRhk8jwRarP2SKiggesbrRTITL00/oAprGI5LUa
kWiheQMsR6Gc0kRznDKPBx/aVvtpzaMC58V+EcRYWSwo0YGrvrCqcYPqh41ilM+D
syi3BQQXQQ/4HTTQRHSJISbXsjSBlFQSTf0+OMA1j5TRsLabVCVZQWRuWd6yuX3n
Tsz50ajxbHcA/c152CIRjIJgbiB9obaFySPsYmy2bdRdZC2WAUEejHMWpHrBKC06
J4ArIvFDpjApN9lFnUqk5jNE+zufjHQ7dj/8exRR8uAkpmtrLKC+zs0QTIdamhKl
CXc+f/t5iBix68bnyY0cdWk8A7hszXukDGlmpLpugOBaK9T3BmLmPr8D/pG0mzpM
Y5B7v+UB/QzxcP10h9oBXzOrWqwQGlGXJu/afuaC1XFzI+ddIduFQZIuUwGvO452
sRBZYp1LVkWL5nXVDuVZDNYWm2TS3btKc5izIkJgLMZSuClIUbOyW1zUEnIkAUKR
TffHZSKN0w54SU6mRpHdEXwacPo6gfbylmo0ZQ6Dx+pOL4zqEAXFBLVtCpG4hVmx
9djqsKWNl/zPF3eT0atSg81/Y1RNOChzcvZxbxzjWKvd/28KZRe+0GgFtTXadDpl
Cvg5jIIqVNNNzzbR2FOmZX898U/05WjAgM6eDpfn6wCzyz7r/Z8isrogx4D6zeVW
xmNcqVs5FokzR3mCgRNuv4HKet0BkiMPXgNsmDgvw+gXRXvaZfKaoNtk+Y3OH3jM
Vv7iklfKAtNtIYFwE9GmFDQkGQxx2Iij8j27JF/njF23jolxF1xRz2jivU+Ltu6u
mGGTFmfqCeO4hPXjqufbVikZ7svdpMzcIVYO5eMaDx50paA1Lx48soyT2NwYR9Vg
vaj9fpSC7ZA4kgGXrbXGyJI5xHeGMw89kXySLjyjL73JjS9G6EFGhdkKAhRRMyPo
e4TAmZKzL2xQwlVQtPQ7IMiCwNsL0NrS9gZmJQWY8bd1hTKXRMXOuvjP+aGE+gu6
rlbvf/+d0v/jibaGEcrLizZmqE89ImZJolkXi/XrY4RIUtaHhJIcIwrlntUIz/HG
J2tkY7qDpR6sNn4E+YrFqkblZBDCyaYBpHwZPvHD5bh3b68Xj727lHL8CpNU2gCn
VOiRv6mq9+GSD3AZ7ddCIzf96FB8+LcYmwS2tZcBSVUNoc9y19xuNdIXMYf+tZRe
YpQACNV7ng60awYnV0ND6qHbFoCPFSEQS3F/0cXXPDmts+LxRlLt3uLcqrT2XzIL
To6vbE/uyVY05lpyi8Gy+KGAdXmHy4mpXzO9b4BVQW0hvmAB5cvth1HSOyXjhKT0
/B3uUlYZsGoVHyGZSwy1V8xYH2s4ovsTGS8hPMw2MNN/WNboB7RfavyHHVTDkz9I
Hg6j0UVz27wnhyxiGDx2bfDG5y3TWy7UeTq2rjzzeZkiXIeJEq18BmbjGn2F0I31
2F6XWbR9eu8gG/CHrQLw52ozA2DGeRctJWz+v17QFAhCLj04ARisaMsO99kaB0DE
uSXzBtzWfX5GideO0Str/inNsSwbi5wLl4+sXzay2Ub246JhZDXHSVStqcUODrS9
Ioild/I6BgWFAel4vSMwi8Dv6c+IjfKwfhfV0YHRqkoIjg+F7Qwm6GBArsvOkArQ
4PhY2xHqVhnMK/9cyOLxIKSQlSG5ZIbt0IDJM87ZmTJZizDKM9H10wUb7mDL8XeH
MNlcJqbfqy13xJJyidEiDvHoroY2/SxLBoScvK//OCJuaRk87a3poVO6rcadV3nF
huj0WHLmICUGlh5WxTXzX4mItug7ykFWIn0gdbqUgGmPfeiX4oukU1bCGxvOzs3a
p7vAg9ZpnC3KYNwC/a6W1k9TwHFmIB8Rzxo7AUcddMCoCf16mk6aMg2ghzQ3Z1oL
rJn5vZ2qp2SW1NcbqcSsm8VVEmxnMbTJlzEyc4OadSUaLVM50F8pvWAvkDKLe8YG
OLWaL02Vi5wYx/ERTKPp0zsfBisUveDPL+5qp+dnmmtOmpor8j4CcT7Yy6lWOkLj
gcNszNJFuu2ZPOqlFtGGUZz380WVc+GO5ZoVEGXtu/F6D17h2F8dwkuvlF3UWBhd
gremA+BZTbgGiWaXb579cjb9CXdVaEHKUph7QL1NWzwHXVDQFFa0bZ+Fa3nHR//y
JPGA0srklryhLi+3NFd6zAe3lbvqG6gBQDvcPNvy4AA2kQ+oJxMQ5fP/jja8KOzZ
HD6i2AJLrunqXTLBM683B94XZ3UkijluYo4oOyBiIk0+dtgFppI7ZWaV2G04hm36
N0VY03+9egucsuNEqZFKqfgpoqz7o9i9q+gH01GSpu6gRkn1+WnEXQkpnQC2F/IB
9I5Nx1iFIUVguRDLcCGsyJDvrZYGLj1R4t6GlCNZx31A6Q2iRcenlFpfu8n1LE0x
WC6nLMOqUQxIbDEvM0gDruc+lUR2NPPaok2Wp0AyEtnPfV9gp2QB4A64h6YAeuGd
1TSRK8WnEsdj5q/V/qxTwKRmKjaMOVcx4Y0Adm+MjIaZRK/C0JgvMS5LSn5myxF4
dSbupKh6qBpi+vEdxtF3665VP8FUVMfV4BX0rpic3u2BXm8ms0qVsEhhX0SydLtO
forGOdkwIN+91ZXl0tPIksrd+oZ21Srk9cmL0VdRaytfkQGOcv11vpJgo0tGnwOJ
cIVBQh88XS2Kw67KaHVoPDrg/Xu/sRnjQsRkVh5PgpLp5EOetsaHDCqfl66hXWEw
Z2duGOeIU2Pmi0s5L4Kx+k3Z2bgXZ2k+AtiiyCwCXjQNO3fWc4o/ji5/svjYOV1u
JesvuXpOZttvCc2hiqc4t6rtxlUA9n5e0hodZEmGnDzhm1TOZj8keSoHoS8uglfO
JaLGG54WNBbDwpkd196sKItJoZVNAr0X8baUUBJoQeh+VBYdDaOW3Jjk/io3YWTK
0Yndw2zjCkQ9yiZiomV/t9Ev/i3HOFr7CQ1KV0SqwVu8SreDiJl7QJtYlMzMnAQU
xfpmKyw9CT0PYAxoLZtv/besw36f67+MWsC3Hue+DHedDK1L15Zirla7BQZp/Vhk
glCNjw5U6fMfSAoM3F5ndhhssEXfIUj8AtPd71F0TnU/Febn6WADZjVomMQP6RJ/
Baydi7O2i7k+wQBKlgW+1VuuBNWdmwcbJRyTi9U7XVLC43Y52uiwO8a45DH7Nqdu
lsIbjfoZkU7ZcCIkQqE3yxkUm/wgSdquC7hHlF5K/Csc8t7ijaiZyDgn5Yi5b6NO
ag4vLwYKlQA3pFwCF1PczVyxslw7mq4SmPAx+0nFDF/rO5FfKqi6m/h3QAq/gyG4
cgKtWeoNSKfp95FbFChhEFVRaOjJaSfQM819j3Jb7vRjW2jaD3jQFKFCGaPhAX5z
1y1Sxp23AP4BXfLuJ93Z+WQgqCxkucfS3HfQQZSjWjBigpFo2Ae9F1tM1I1momRf
aIeIa28fBHQwX69bOv8knHrsJCO888wOzJi1A6iOzyEo3sBl+bE9woksGc+nRhBG
eairHCRX2ebWaGk/vt0yUDcb5GuMjhKntgwahqb6+wrhuSVUVCOLobdgeQsDIu96
LffBYSDUT4hwtBLWhhV82Unv3Zlo9l3x8mdzztkfwc7Zz6NwSX8UpPvT9m1SA6SQ
upGDYrddk7Y0ktyotekhjgY0bgqKjtZwThQMrLTvltp5NojRD57BBkAT9WRQf4qA
9z7gsHqd2/mTl3pDucu6YGyOnxuJzvfCmyv+JtCJMXqE8XZ21B5R7CrihJl+0zHs
9eIAyldnyqkOcZQwddO1dY6RFh1hEbxzVZ3Sf1zRbonob7digXL4DVndsViompgF
W6iR4s3RvhNkzY+xNKm4pGsjpCfDkew602FLpzDHWeHb08gaJViZAYXmNs9fNwgK
2q7fn7lwKQfLJLszNOGHZInMOOHh605UB6qC0wzj11sUlY1vu7/G3ZICrxGu2Wis
znAoPmRg66nNeHMJCvQSDBtuW8L2rvIZZqOC8CMZZB9sw+zpiGpdZaW0PTfJXD02
4+f8v+U2LLN1E82LZ7sLrUmRopLk/ggOK/jo+lp6W1qHPx0CFBQz3UgiouiGRpqU
dXW2k79EOnamcy6NlQa3t0X2Qou2avcKKy297p4pgaqZMGxtYKAlqc88t/2fJiU3
ZkUsWpqCGSFyWiHxauNrAiBAXwBMUlxIsdmyKnl9AHd0gjUVGE5I2Kc8xdRPKf92
WBet/5Y2h64XjhydopW3CXebxG/huQwmIQ8UGiBkl3XTOWL/0Z/lgMbqgftnapAf
py5qWa4y1ztyhC4T2vzT49Sic+hQdt5oKA4PZklG1bw+KmCxCrh4oniT8pDj4QsS
rzJ6TGE2hWWsSefgrA4lv3S2dJgsUyiQCqDbp71CWdVragDwXYNo0sVnia7pAzgr
1Vw2G60BhqxR1alHWJ6vrZipZcr935s98NJj1E9FuyCY7GfO66KIMurYo4oaC+w5
REGLRa5N7bohtj8BdNhgwKZrTKs3OXvrIa04LO7b8HUm2lJ5sLQW0Qqh9InyNBwU
ysNTkhHxTELZ/VuD7YOcTl/JPhQIASaYadYI4fI7F5c74Ij098B+fFqCnP+lUXtT
PBD5jbfi4oWewmo1fdHaYBUvZrVY0rgCjgKPRAKvYWVgX+AOOVyoxOp2rhw+N2AC
WpmydAhPCLpkAU30+8Afrb5ouU1KjLORPNTdrTKhzVlZRm3S2n7TKfMdI/nVsN9N
/vkxOT+nr4368F5J34Bqjtoj166iOr41KF4g2ERt4PCmoMXxkeTQtBHcHk+UO/ml
YuaeNSlWeJMUZ9BxWEFxK7demFRGs0mtrbHC/rEKrN/x+skvBa8WUhAZGYqSkDJS
qhnbkNmCFW5GaWExWTwNWQM2tc9hUjwgTx1jracEjHrE13XGTOmqHJSIVkxT7GRI
oM+tHgqVpRXKGqzq3SGf8VyCPb0YiSv918PexvbDF5nhlB6chHu8M1Tyjn53zv5j
WzXei8rk6o1xnVtfSTBbUqb+yqAWnnYHOsFrKdP1JnRTJ4I46dLSJ/2d3iYrx8n6
bE/gtNs64hnnjFaJqF/tErZrGTqJOtVSTBg6Tfc3cATrnm+mKzXwJCX1sKP+8cky
T3761XQr+dZJ2RPriH8v9ZG7h+NOlrBUUttxkvGbIT9xAh8AUkjS7Oqk9phclEuv
Z4t8wyfDqj4u/zOoSXWohwrLyx3OhwQZ+eGbERmQEhaOfGua2P9gQtHuV3eRcMif
wUKu1OBUIfX6dPQpmRlsrhXwVh4ZfRhupTFAqOcLW3bJFIlwWrHg+oP46iARuGdS
4jzw9yAHaSVG/n8QOcUt0lOhjjmw7YJasZCwjiXGVe5OXWwXxHGTF/aFPIc3eZFk
2iySEYi8TYH+ZQmuaECT9VHzzCxQe6Kx7D2HJ+9wdPaTgkuokJ7YENPxhYIavfUz
r2VZn8cVn/a2Dr3uikFY1bWi6jiiRgA878czUCHuxlEyHbAB9FbIwAGXAe8oj2U3
jwbZcVSPz3ITf1e6bQFLDfPd7e7xyg6QJ2jSV2PJ3e77eeamLNUqOS+Qx1IL9TMj
iWPzErmMEZKMr6LTkVbEmp6diX4YsYjyhhy5ARYpz0peHMZjzFe47uCGOwPXvJMI
GH3VGgXoU+Q3XjZ3I1fBwFQ45LQaJHLO/QbCmjNaSsU/4BhsCbmy3Q5CgFs4UYAl
f/t48qqHXlqqclJ99Vjo6nA8pMHzXqZL7o86ZTXvhyCg/CYdkKLzjgLa3B1noMcy
Dl/lHgfQ0HNgLDixDfjKSC+IWqDboewgcBAutcYqCoKxSNYMiAwR4uWZXEULPxbY
XVnnX33Wq/y3ZwI1vZ/XSB1mi/DwJwLTnNPUArbltv0yNFwN3pf6+oiFcHF9V9OG
8F2avmzJneYam6fwnt/95vEfeD1Kgq49H4Vzo+anEGAI+1Zjqai7te2tP7g+odHC
Dcl9+eqSbfbgSezZhYpV8xUyUfuLWnK20MEDqsDpY3nFNU5JPcB4D4NFdrgi1Ogp
6DtOz1YSLj8Mt5v4/kamxeqOZc0nXC+IepupM4ARvWklye4A2WR8spAOXQnNpgfV
27u/kxyrF2bm/Q86AMPUt8Z50EQg6xzF7O3/Fu9C9NbFIRfE58RoklLIx8jiuCZr
biY7LEJhvbwzatph3CNjVBLN7+AM4pF0XrkJW9jiPhfVL5ARRwO9ZYJav4n74aNL
GUayYYJggoRUmdaEUYIyFeen9ffuIKWIGw948wGFADsX7aiB8Dy8YoqaIOSDGyLa
aJo4B6wN3tZ4PIWyNelOjJKrgulFrQUHANOoENXVv8SyPFL5vUGFAyisWOc1BTFR
0u15ZW3snmQTdYIzOPj+NonTMYkzBeoe40BoElFeB+XUxLiYp1KN3NiL+BPsS7tW
2Sj8tBYCszohhTqx0I2mAnX4KSVD1/q8h+WDoUUNw4DqbAgk4ORf9TiNQIfFde1E
fdNkPcH8DN/TCRIa02JTsIReK9B1skQccWzw6qhrWnMsf/5VPqC6wt/gQVW8lwPx
Zx5v5bN9rbayM1+uocPKk3W3nyMTZYkhbP5/NPXs4BvksbHUKzYi7LqFstdL7ijy
tvCMR1Foj4lMjdAJs5d5g2yZGlw9ATW4E5WvwVitzxObp7f4pDcnpvm3toleh42W
oIGWQ5w4vBR6KGuL+xWE/IJJsq5ohSfUZd1Qs9CmEQJZIKSzJCDgzigruNojfS+B
zdnOg+nTQy3rAowWf7yPpSYCvh33pqtJIBu9ybpoWojSqUWHVyBjey0zUUF5ZqnX
IvW7GhT3+GyWH5i7MyY+UFfDADdO+CmiNYUbm48+0zqauC7L1WihCNfWuBN+Sy7w
1xdLAocXv8Zte5YQFs+gi350aCUeFG6Kk+8KLHq3KgBkrcBGZga5ll6ih+KG51kq
0qopUrbzDJuK1H/qgynKPV+SirK3G8ve2IBFRDpnVCN7b0WChFUwSIprZmAfUYY5
pf+nYorQkX3YCNPFY+gxxk8Gw4IcK5WNIF/5210TWO9pS3OZDKPpC5cb0yiRp2uO
5qxjjkUKjZjfnk+7AYRmBrRU+DGs6G5Sbwr7qOI+SNCLiSj6n1L8cXB0V4l2lanD
kdJeEhytqzq0aa1d4xS5gHcff9MYwvGN4Tl0FseHQKrnxj0VmlONeJJEhJCmLw6Z
TAsRbRLK1BwgK9Z8VdgoIlUu6idTURlOeJ8DTsEQgn728yC1/gF54jdZkQEe5jUl
vZ0XUMRdTOf4DpBaM91cfAGbaQhYWnwFx0R82kKHO/unkQEQlrxrdaEYkEDOLHCL
mBeCXIVnyPY7JgrxncTTlsjCD7O7Oga00wvXafLMqv3roKKoJ4keZWbHZ6rfgbTE
rXq/9fPSi5r0QRbicdh+FYHaihZET/6304etGBjv017/nltJums+/2w7GnyvGZMl
HtPQ/9hFP1KU3crWumupS5vUwiwmQoaDFmcFyewYrlwmz7jg0SjHPnAb9Nk/GKTH
zhqQCB0YwAq67MChmrEy3wHA5PjnOsEQnfn5+Ue2fWd0yGt9CMPo4jofA4X1y+NU
7RXA6sEeLBMH2BZ9ctftEib5AFGX3l3+g84AisSsnXE6W6KjdZI5cKlilBB8x6o/
RPqz0oc8DeR033X2Hnybyt+45agmgZMN2fm558jY7NWw7ddSWC7yBKr77puY++gF
YxmVg/jCKLNZkBtjyZYJNrttaax4qgid3JaYtOmC9HtgR8IhRYJdBqBtGMeH6NYm
Vt9K38+gQsw72r1VBdPzaPVhNUvXtM2hLyKJrtQPtpKqwO3F7J8yiWvElMjIXWQJ
fAldWsPunwkthVUnOmbdjol662CdKndgUmMByuReDhzec9LaSN/oPmNKNgGSmHPb
p7Tu2kI3mH2S1Ps3yiZRse7XIllYYDRozCGDnqNWY3+zuBZNp8ozzqhWMdR6aRrc
59BWkIh4o+AlldGUbVPZrPpbbY0xgtvhQCNZpw/fa9FfMczsYibRbIRQLLjMLg40
/+//xA1wKv9gXQvXUi0T47hTOGEQWX61u8awwsS5Lo2il7bXzuBdp5BdK8WblRnL
3y/4mUcNAmZPS4QsvXkVoAfuhqxDImkdwBewfBJsfXRqLjdBwHEor/PgqdPdzIgE
zD1zXlU9is3asUsUbViJ3x5JBrvdJHiwZWBRJvpZZBAPbDdRGBLUQ9SewFTy0Lmr
5fFguFzx4Dyi6lTO85fjq8V1mJ8PL5W6YzzbeaOtsTHwSdXsUIm8g+APSmFIkUeh
sjoST7zkr4XCxYwkZlneK0fDz4FcQ6IWxWV2Wz8iY4e/ja4a9yfjJgeUgGDZP7lI
bD4xE3hC+hFsH/Mzb6KUPVpQSspQNapGIqlTSWWWjguop1n3UTHdZ+hSZpkwAE7J
OtoYL/uou9wQ/Pwn0syvwjo34244TcXTV7cNveA0FZuBOs0xpwUTTqhQ2BnQxLFK
+nW1QSMqbYqLSQx1YBBKonTM8GcyIgu82uR0CQ7U1TrXNl0ZJXfVrYabRLdfgPZ4
shmSEUF3FTiLT+Wg678Z9XMkD+/nCb89HFIM473DNFrrlJMBGHdjHW9X4Ve2SsLz
LDaPdjVqdrbDlsbukWjoddDu9xbq1Ptq6C2HwNajUQTfrXvZOjBs2SCA7acZob9M
83kHBYN9r5Lta8G8QLwoicYmXBAG/ph9HPTuOAtzHQXT+rwImQYKByy6ImRrSAzl
aG2ZWh3HS6jvL3ZZwDIzsxjSLMLLPsAGg08AGDMvmkS4SNHqjeT1PpHAxjh9YAfe
qJpe3pbskSGNY+cDVhPH8lm4DBav4bZKYe8hPZTnSwT++1fAizLGGLa4JKloTXAY
J4hjOAxnlDy7dRfxETT3DO6Qix37bdPpnjYNQ0VITw3XltsvalGQ9nYHD1UYx5C5
sk77iz3Q1cmmYpFb/vlaNQRPQrVeQpdzE3kuZOO2FV+bqYqrOrmngJd0mcaqMERz
eQl9LiiLBTiB3mLcSdPPyzYQy3c8yGs7E7VhQLgGqFJNyg8RRDPvyE+hS56plWfe
+63c/ohpg15um1ZaehuEXvOxv3EtPiCkFzplYG7zZJ/gAfImKuKdefE8suUTA23m
y3z+iluIfNC6AsksmHtOWENVfWaV4RTnh2HBXABr7wR7igJLcX1wcOjOkxNKzfnt
uHlsgWsOdDSajxCSnM5Bm1AET9TpPI28n5e9SfREju+Q7+7BuHT4M/evnPGVn9jf
wumsRWuuV4bzEvpwT/bA0N32lw6QSK88V/gFCxPdwyfZvyPuzMeomLjE5WzIggFB
fuJGzoBkfJjaabH/WfZIoy0CO2+WvtiIEfPHllHFFF3YxrVJHFI2v2SLgZUnq3Qm
k9tfDGIanpWsejV0qiaJgkLJPHwT6OCy1GE7COxU9Z+gaOOuD+UWYMn2FZYHKeDR
GFtxlite/GHbQNQ0TpZ70un2v5/mFYroagD31R96gydo2rxGP9z4b7YSU8xNbTJ1
1Cy/qegI1DSbqyYgVpviU4STjwYPbjOzkdJGOh+TXOQkfLwPSGL+PzDqwMgN3zHZ
9nvMo9MaTE7ILmS44BVUnej7JFGZU4GFYFUxxr8rXyeNkshwIiF5LhFnTazt8HcX
5caDOFHGGscukeTaxAaTjlvlGJvzFMhp7HqRfHiFEJR/Rh2yXkJCqUgWTCaPW+38
2xjBGprgMzlYcO7AGFjawt9gAdpva4dxq3GjvF+xoaZ92Zex6gQIF7zZrRBRDlni
sVTurhZc/6D32TCWhh9O26zUV0dXfFnd/1Mp4C3e2wObWJVdYzlu2bUk3+DQzFsn
JY5yQUOJfc/Mfm8/dwF1Zg+4PqlOUubh3tHnFVuFDpP/OIxJgPMSIaYVbSh+6rpX
3mtjejdwDDQynHlIKrZFvakcdP9IAX47HnHXFdc11NSg6OTK3sNX41mvUgaYTX16
n/iVtPOLJ9MBkF3QDKkBpyu/JhASP5ogACR0IJaL7hD5zKXUTkIllv2mPZj3Ep0Z
v7W62Vx7UB/ZeDsqmQqimnTwqEqPF2ZvEbnwYFH+xdS0qqazhm2Tx/H6goLdPeDZ
tXMj4s4OlgBhN9/3Xh2yhge6lYFMi0YtoDWERx0008NI6MKQkyIP47h8IM0KgzaP
G5vdrnM7hfjpm+RKdF4wWcDr0mHk7wa8pTCOTX0xjFyd+JOQcBwQzTkEINvUquCK
eevbv7NShLI93GhsqJErHNS71RIcgTvPmlrMDY0HssBz1rF/aNIFAsxE3V3oZNKY
8xrx4V+e65E6KweEyJCfvtbuq4HkUbVjgmJ3Om42lNTnKZN2LKihk8Tj79P/KEGJ
igry7c69UgpvFkJ0KTaCYRE4D0h/qNlKf6IMcLlYinQnyMeH2gXZ5UeIO88cjXSy
p3vIlgGMCvtxQSvYL8xm1KNhP8Ii67ru5i0Sx2BPgbSBR1ATYsxx1wzyirfRbI8K
Tc4dQKiXykckAta/qgDRD96DGji3Qx124cyYF2kw9MlR94Y7rR3iJGKNrN3auxxY
+idP9X+CBmjLlNVovTTVZBi70JwtJxVVI2EV4jJpGtPT0XBjlUzNyWiPrIveCQQf
KuxxxFlEV6S0tckuGE3i2vdwQ8UeQe1Ylm3V5aPULIyVVnzCsCSD9Fu4knKLI4Vl
6YRf2z6EyDHTA6x+aiPI5FcMZ1WVotVbY+oc5WFBCx6k7LKKVNBFJIWSN4jPSReF
m/ETDleDf3IkWLFijSMawu96+0aw+stwzrzbMGnNbJzbDHic9onttj3VNbbhGkil
05LTZNDiV4iDqv0/CwQT87ThDE68eFZnxDUNZKAWEuyjNw3nUkXGP1P7SD3ODr/v
VX+KSunSRpVb7kBdTTZEZEhOVk/p57NXUYte78uyzChUdeeYKTprayZYgrGT4fFY
BFsEyWX6AnHDE/nrHUGuXTR5WKDNCPqoThJ61fnlbl5cB4K4M92Pv8BOpHC0Fkc3
mLRdS47f4YW6ra5MxrIuIxv+8d7ahE18vshnjPl7aB2tBzRyemtFZDIw/oQvFOn0
PpCRn2XkogYXAGMGe/BN8Y5zoSaFDt2Ejbqp5VCtLrC8xGGs9qIjM97msZc+FVz3
X3YnkijC4RMFYiZN0vZPZ1Krt5nAMm38X2dXIYZZr1wM36btoQH+Zubd7iOmldK2
2ncUGbehzf3VFAPAxRZ7tQG/k4661Y1EPoOOVY0OPbaBNWXuCPwBX/elmpn5zGTG
SEX8nrTs6YW98W1xkvrugTG/VL0BxaKan7MvbPKmb/XkmpAJV3GipELKa77iOArS
8JZz5ZNd8QD6FhCvTbLPT9UlRSYVOadL6SZFJY5mW66l/JgKBOoajhDWqTE9DsZw
hmSZVxhsDnuSTE6JMpZ9ZlbyVEyLKzUEhpSj6nnmfpn0MNiAwQu8IBDIvAk4dIfj
Ta8UTpi2ATytnh3HTy2kGyp+scq2PDpmqCOHfGw0J5pTjVygeCd06RnrxDyWL71A
BDbJ/iiX51lGmB+uyx1TTu8Kar5mLziiNTxe0O33EsnmIfF8NnqNmXL28O7ARwoU
3r9By+9Pf9YESWXx6HdXpr/sUp3FEcNQ682GOOmqjTaqOPaIKWOxHLAsTasomcdf
jDgs+A+Vumefs9eoQCGpJRTWtBBuInazvwSqdlLgAL1TYJC1wJWHx63hVhiHcslH
2a6Pq4Lq7iwsi+VmNbFiVjFh59BtUtMRUsAUXVgIdrrndKGjUEZuugXhTRY8KLU2
mPxIXhyeQVzaEQtYD7P8wr/VOH4cr2HZmVpvnPnSE5OESdFrElEOB9BM0JXzVw3N
sIecC/lrrN9kBFzquM+DwN2ZjHbJf54v9IS0l3zFGRJEUsHANrxOaTRHGpdoRkp2
vp5So94w/aM6ZGHRO61YU9ET4hSbkF82pGtC10ePC2N++jfMklwN4l7+SpgeOYAp
5+bLWHNHWJLoTj9glWIs+MohaPA9SzV4+bZgPTKes+eDLvJmEQIgfQSktUtNbhuc
pe2KywoaNKy9z0w9fSp2K4s8Veg+x9ysVv0SszhjAWQHizYtwa97j4wmN5ZqiXAl
a8dh5TaoEoSLEy4vUMPOusLfgoIedw8bqVMX2CnRRy2E+7vgfMn/IAhlSUL1/7KB
QUSBOCdEXLWrZzHq8ijtXO+MCIGV5GRJXhlTPY6Hwlped606u0IUVGXxWmAXVBy7
yhBafgQczMVSFGp87TMO6rqJG949So+iT/iA2UUH+8TUHgFr2uL0ZoV/vUTpYT6K
BuLbZH5zwQV/5rlPN4qLGpXXIG6JvKxbJEAu6ROu/cFh0ywIcgoGn9VqKRsAyOtk
948l/kGY4pmhGrbh3dVj/HgfqskjUASNbV0UsMvF2+1g/3JNYfie/IIeRYcmXaL9
mwXdPiQId6mUrVvWOOC4alALgFBUvHI4AO1ar7Kex/+dBfN+rC4GmObuDIZorrfd
cTRLJ1uLNupOu9R+69w4LDx9GSJJztUqx2BEDA3Nkw6YftXawpkdKJUnWJQdxUK5
yQDenjyvrujtyj9AZ9KK8ZZd6xx9gsubwVPxzLIAVwCM8vonjWwWa1YoJ+wh6yIp
j9gma2uKZRr4QRd2sc/99RG3oNWZNUxBJrYqZBt2h4ZEUt4q8CT/EBV9rqoy7XpX
+bSpOaG6qAWS6RWAqzH9fBVw53RSDHfDoJN6ZUb2Zfjz7qWKE7pMKLZ+qZtzc0Hn
Flfw5pV+RDB2xFLaCsbm1ku7VKpgZYJ40v85wl8rzTvEMkKZ3Eb0DkLbvVAskSLv
ecZ4GBTGIhBfM4n2AD2Z/DOxzaSa6R/lQMRRVl85evMy2gnwGWj4x2J93MkNu4Xq
VrBGVahP3BbQhVD66U39rUQjwAMtq4THTiiDUZYSamhf5bSelEQkRJY9C/CXPZvZ
ckPHcmhxD8Bc/x9djB7cF3eTmJkTTCtJ/R6iT9u/3/5qiuM/gsru5IQTTuD+I4hh
b2nHo+eNLzdorEhsiYwiPGP0pMYZDAfAE0GbVAT9+colhXfn+e2t7TQZ2GTsdqm8
8M7tIG0CaZE7WWXxdvzrYfgEvHfagnFjgI4XlFx6/1AmvTLRQMFRpyBL9MoclE9Z
Rav0/LkMUSFiDhBkWE96FpFK/As9ITCjRAuO3BU2llqGbadzSw865RfW3tTEozBV
3S6Z6+4enMacy2/TMHwp7gzIqKBBy13/5tHaZVuCrAghmnHzDQkcux+cnKCWclt5
yJTM4vuzJkmURZzDGPNQJBj0CWGVaDXCKtGp6XvQP0zLnennU0Qhak5bE+BL5/nf
Y4+lTWtlin6sWfZarWlk0kAdqJ+QrAV3GhjLAWz7GrYs2wAuY0KDqr/XBTceBTnS
4hwt4/qMzUWgbvpir3gTwxu4r+f2H0ajl7Qz0zL9n2Ev6M+C0MNuYpEZjWDmLIla
UyoIpyqPxDjb5UO0ocdaIeh43xPBXRmxuTcmJEK21rNW2mxpi55D1To22gp12W5z
XlEVSuyNrmAeFnCy8zfFYjtc6aCI7qVNRW/YrtIGG9SSnzZL6V5lwWX2CnJqz+it
w8covtFcvATSStsghzZApUUFndD/nVnBEC+JrkBmcBxNDkdyhkKhvPKbc+oHErEW
BM+hHerNVqEjvf91r+kDjxeK+jYTnKsFjloh/w0jjqLi/R1b/xewyTCkk2zbqy3v
lE0MpIUE5XhyRMf/O8t4fpuMN2eMFgaun06z6e/v5nCj4H8LZ7RFeHiP30DkkS/c
iha8BqXczcu/mDgeXMZjCRhKNeCGGzs7K6OcStIdLqAR80dQQijNf6EQ39XUnrHQ
ogzBLibOiPca2r5C8ntTc0REF/Yw5H59Lq0gPgKuF5PY4/Iqzf4AXQw4mmMTmt0Y
ZJzwhWZviK5cPE0/+eda4cVe4nbnEpmZTv9c7THfm0W92JrkQjQuLkD2lE0Sv0Cq
wlS62tJr+/fFoGU/KGWJPBRLvFu3EQYAkUvm4BL7gI3YwkmvT4HHeUYQ+mgM492u
EaqBPFJ76kt6sakn+lebUvz7t4M0X1Nh4sSeWglLPOgYOLC3cp6Kd8oBaKwG2Hy1
TlfBeI/67bL9Q0qspQAW5grm2X/bZZYfj+CPny95aSY3LOJT8VLW0M9s/p11y6Di
qUJHaSdjGjKxM6K3644xU2/r6YXgGVk/yU63HLrEgS8TCad4PatwsJGk9ePBW2ZC
Wl4Lo3hbeC0E6DlCko1GqCWckOEJY5g049ZGZlgF+Gm/KRr6DAx92FEeq/ZuoK7C
klrzC+1g+5IKGC7e9rW96xgwnJA62RzfnvV+4Mx605ClxBKFzwK94gW0iUvpbl2R
+eqU8vgAID/Ng023S0GzXbl92hxgPTJPh1LKjW+KFsIv2YBykGvmAgum9peLcSqR
F6NcmxYFV/KLfq/DAt4irbGI53uwwNBS2T4UnZrROLZz+TNTNe+g4y/4befpsTRB
fthNqWzIIL+/10ZEGEG/32RajB14MNsRmG6IEHwAG3vdUUiwRLo3cjO3MBR3+oko
nLPJf/OTk209pFVu9Q9RNKx49QzTdEaeoKfeRIwiy7k/FL+X2+DWyBCbukI7gJad
LoP093Fw8JlZca+hzgfbnate+Hn6K6kcrsl7hKWvoeQxPTCArv1GIIaeGtVzX6XX
v+T3vA1qO5zTUrfJAEPhA59NmosW5WnnEetTDeaBFmaWd9qZCytfYJ5puQqrnn/I
J5N/K4AxNzRavPlwnJ3P36oKwssON2yeLL9BaD8hF33dMum61J2QeTYMForp17UN
1HHfiQEqiHpX29DQIpI9LI6bcVdd289Wwwz3Qx9JofhqmsIeNmd1erpjXIRwiKIZ
gKL9m4+YdAY1WVRe9EJ+mNdhZHXMmZ9DxvEkR1/e08YRtx1XU8fGlF447D7mvoXJ
DiyvKHLy0ILk7w87pbE84mqKxfjBTLUZ+IJFpIBy2pM+Q4BnHBxkKO58CKGc02gC
WbABHulrD83kfJgJaIfr9ddmdL//DuqLQMD+150lBVRYnisW8QcMqJj2VF1CTQht
cZuDHqYXGg0RpFcJl9AYFhcr5t47iR4PePdX+aG3VVXippV1/p3Iik2ezcgoNG/7
wkhizxTa/2+28nvC+8V/v0JlYbe871wUG43CXoTaCqeHdIERNIU5Vlz2udpdFKSg
IoVhI02eK6ff92y7Lufpzykd1yIOKvN0LszjMNYE7EE8iJZ27OCuYhjsdL2YfsPC
ooxqQk9UEpzgOdscR0sgoZYMUEsMAgerJdsRq6F9NbyTIm/TS2RJXE6k13LAnluf
iUpH2QacqjxSWrKE+C8P/avXGE/Tm4pw6T+STK4I37s+stEWNljU8SjCnWWdvVLG
iwOwdLDlrIssxqEmL0GWU5Rys6DTiU1YNzeU8by5B7Mr2vp34jS/1/v8FlGFd9Fa
erbsh11c/caJOBNmpTw7o0wOW3O9Pla7O5fhV9/+vVPi/Diz941LfohQjJ4EOlG6
fPaFJSkjylSBTcxLK5ynAP1R93nR/Nu/XeAw3dx+mrWSFfrUMWynk04+Y4xXqB7B
MUSp7VIYRUtZSfUqze3ZLXkDxYzs1ny4W4Y3ozZsUqCndmF0z+BkXAnfkcBCzIcf
vIJ4YVAe3fq8X601SXgvOwuf2e/6BCSuTBbmTkOOZbfkBeEEXOBdG2pB7ApwSRGo
X55IBpBYB6ZrdnXlRQo8cTZMx/nbBs+X+zGVdiJ2ZH/kt+UgNRkvjvjCsJPLz/Pz
qCKc2zPNzjBFLYQ6Mh5dPqQ0gEZX8uP88nzmSW249rf4+Df81gkjbVPEeNs0XeDd
0Zo7Th4t34KBkbhwCDvCn3OaZUrWjY7gRxhtlAkjATvfDYvFTkiwO8Eh3mRNMHaO
otpTg/IANxJTx9gOWYPv7z5YrBbKjwT5KW+uxOSB4ZyigsB8hp2jBZQjHKIcTukw
gp6r6YGrs77y0Pnrbg80Ds7e3ooZrAe4hOZuxk/v4eogV1jpFbI0rs434pjnmnX4
RDSd7ADHK+8w6mwtPstvv/t68Ke2qunL6Y1GrBp+pe8SIstHie/8PNuSsmNucpsr
W3GGVQTknwAAq9sfWBoysQO551apDCnYkHa3i9MRkPHWNpoAovSPJFD5Hd+Xaoej
q0NT4GXLccsv51lf61FhJt3/t2i5wrZZaVsUbb0mdoAfmvUhuwP705QqLYGbWYed
GvWpy1hYxLpoA5QH/8NLE2fiJkNoB9JkG6xu8dva9ehKHjAPWdV0Dr6VCkepPFPn
lUCDqx8IDGfeNiuOGlSTP0zx9BMY7YCXgpxSkegZa742SeibpOFDug3/F/OLA85D
e4LrwNziLAFbrYTkqqcKuHTlB1p5mwTAZZ2yC64KdtYE51SG0WER7WEMmgzY5agc
JyWP2m0UTM1uKStdbrwtzWdgW8bQfk9NcEm2V7N3VLq7nuZsl3j/VFIStAz5UtnH
sWE4wPU8iCh+5FpeCFNSbiqRbLrDjtpqpgr8nnOlka6e+B/YWQFjbazVGPBgu8iO
xhk3HklWIJl+9t68npWvC5/hqMhx8/zx7MAcsOt2XDMozDdaDXnZcihxjWjd+gJY
KP4rmffHQi/TEOmcBhfx91yxX120m8AV9U//bCFJbXTf2f3m695yuU65jqxeIyJ4
0xxUhuqmuvFyU35wD1RHTk7mwHfsPC4BGHx5BB77RKuUBzsslRYhJtXEIUlrd7K1
SdQRgZV6Lk8FQOV9J1FxEs1Eov/0YFLm3fgfdxCbHGIJCSVZaU4v33r02+lapv/1
4jQpkPxwh9u9rhAOFH+EZe+eNyTeF1F7AAL7uXYf+vP5qo+3s6kXssXUblXuklW0
QYnL9probE9zrEoYvcT84+sSIqhsp7BnXg3GDikwzOQBQbO/A5ugLmOF70L/hLc3
bZFuGr8MxnKSHdYLVSoljHN4H5pOWluHzAQJgUzGcG+TEXFoixQ9Q+g9YUaeqNGN
BcVYNTdCiaIxFGb6jhs+uYIJOqTKL5u2e1CtCoTFV66DJwfAQmkhod8HFh9vzLlD
FxIQN6XbHJUKNhLCA7fg2/URVi3ZaYgsmL+sT0Pp6aOMHdx0ti4zZrSyYHYh9kJ/
L0AMGj8858h9l9OGOIbrTFX6Yh73MSZfLppGdkVkKguLYvGasvQbneSBeIExUaAu
UHeaGriHNH/+aIH6z15nbWFMEALTE3p4kEMqj2fiFtlXwrodRjcenveBTFUpwG0N
bH4UxpCdOEsXfjCyI6dYntfsTaAi2Fi0Lm4dthaNDQaROVAgWMatNwvMS8qo0u/V
WNWa3SDYjVebswRAJA/oq/Kpv8QbFHynmCUrFes+W5lyPNqus4cAq2nWA8tY5SDw
yPqzRsJD76MTwEvthJvQZ/LrmKuHzJ1tASXvd0U8KTyS8w1ov+Jc+ffDOGidO6K0
AeyCy1XW1ylwH/6DnmcX5aXZjH2bWOEIOVMG2kob1XisrbVHQRp6nCi8GgAopQOE
sfBJWUggiLRIYnQOOr6uTqbul22nJFUq332VZQUamgJ2J4Urx/I2/6zo6TvKRDXm
2yEHxEKJwWTFv072M8HsKKDIxRhUDuLuMJ5rAE6kzxIgBapgyAwM1akzfrXQgG4j
xFQ/17G9MnQewFpsSeU2MUe6Kk2DiPojumRdRL0uz/rE6WwpYzq0yDkDzK+uQaqC
Y6GbHd83mL3GCWilREpSfMFe4jtIZNykDRaiPABRYfRJFdVKqTpYrMg0IFsRbxFy
g/tndgcCyP8u7+C5uG3/+VjBiyr6hUAtMjPwcWOhUiaFwIfLMjpX5hBkAJW6QXYM
4icq+NVyqmkZ49c7Roh3M4c3ngWTHb2ivh1Ljl+zuFnrkfEKsbnJYI2izZtjfHva
piFdBzJMmlrhe7j45mgRUwDHJU/WNfkmiDhvNVa7oMfjRfdTo7kYPBXt9E9IR/Yt
m82nbNCjCu7bS+TkRH8QAp+D3Qq5zy5ywGFLy5Od5eU74LyH7B2GErn02lYr6rcj
RMZJjHV28oNpZ1M+wLrP2fHTZRydgi3zR/g8HlrqGDNxaKHVJmJf7w3GXyCvctN5
rbGEBIU1mGWq+atw43gnq7E5VMAgdZ5rW4bpoxqe7qPaDKqdbUCx6MLTM0fLzID8
R3rK4yhVkqQx5hXxza+GoSJxEjVRuEoQBaNMh99t9TSdZ7d/Nz4utyMChROFDMEz
Rysbh9tDnmoRKZycKFL76nFtW7F1RizO4Ur0iXj196lrWsvsG2/dF4gaeE+jTBeH
ASTw7+Rek+eM5biMJ22U7iRSqZ6C7M0mRKPyKNcKB1BT88vXno9yCeh0afp2e8Ed
MoywDJ75VBgMTUJs0Ysib7dddA5lhSYXL/3F5MtxpZaPuU3BovE+yDF8Zy/lT5tb
tcL7XN99GvkYU8Otp4S1/oS5S5UV0im1RxPbUj37/6mTPWYO6Mcpyvm+uXyJtrMn
UPBIPA1Z1uD/Bj+V76WiLgJ/vP/tTgOwzpHcIXgbqizQPQ1ipdCZc2kz6xuPsSNI
0+fZPQchZzu7s6lEOJSNsvOXv1wb0XEUO0jS9mxuA2u+m+oSFHiTYv596DCNi4yb
0a71WA1fUTmChFcgEwnOIhF0aeCtN+vcuQm06QrRHxf+ci2GG/Xg5IdR/Wdk1TNj
GaJcNVl0scC28NotPrtGSEeTgnzLQ6zFcKy4mh9nSLWqSm00OgWYHARORvx8yPwD
rfJqMKywFhFmxPLzjPFrQCdhwVq2uXbXSD1CWPAF73fWP36xRs/1guUX++NzEXTb
+oCvoIrBSc15WIyvfby4U9l7MoZRw6H1t2gPucvPgxIvT/VfHO8CQLh1C3isJ1eu
VgZI2hoWGpbrWDhKNkwPG3RtmTpY196JeKEd7x6PsBoU1fTHFjO/P023w3iBduRK
ejacVxwmgolqtskvmpJIMhreehHf/DhsJLjW22iuvObMhlBJ+UmTW1bLXHz14ArK
gxsJvUt9K+q90pg85MfTF+THW6ZWjzXhGkFgcAtelnYckwWsmXmZS/OhsCWFpw1K
/bymdaWnRg3Y0qLtGmDbjPqmfx+e2VDPonwzE30QUvbwdrBDZd/V/2UguON1q+03
28t7IL6b7uIkpnI7HGg0f/X3b944IQAiYOTVs4Upx3viDmQoi4RS9AfjzN2khKBG
iHeEg8gFLMHXEODCW5GzPX7wPiqHXArR9+D88Y4FD8jU/cI9notAPcAD5O15PMYn
t8OPv6AuHIpM740xGo4GvDOXvJNTiinfpIb72m0z71C6KuQAMxwoTygp8af3/H4w
GG79RHnC+ChFTJqfCHIwVx/f5GRA2ItMil2vL6kmvHOnZwUgIGh2cD44d/5Y5cce
qa03Wo4QfXbCCxgE0j5nKJBWmVTeyVKgIkAkPCr8ROQ6MHf27DP2VzoQzRDz0UJL
5Jz+a58V7PMzRSPGgXWZiJKYyBKuz3M4rwJvxadJOuw1+uEeg1GUV7N5tR6FW/D0
Rz63RfnbnnWWMaaL02Oa/w/MiWYriprRX9y90ofixzpRGWGM73inrVXaFjB6T5So
xqyJxvF12zgC2sXetQNfrSk6vPCbOyqgs+ud7g3555wclEDWfxblx+c66gUtzDQt
Syx6UKQDm1uwAWOTNnMBnV6gljMIzKyDloOXoTNFAYemrF7aqyo/FcAZELo6690L
b50X3FZnswrG2F1TcQIzRLEmvdcf5/liIp+OLjnLH2N24QrNEbF1tszpXsYuA6Hf
agnzoEcJ1ENkvs67zKTXiDLjzGxXWhiYt6iH0n00aQipBpkaEhyE8zSY2HSCnnup
/X7ceVlX3UEuZ//2mom8bQTuSjnu/iVdTgV9YjkRp6VYQ4FA2kgREOfPrEXVEXEz
98CgPTGeDLstNAt/d8w6+HQFngDBCa2+geKioKDHC9fA5MjgHtk1TL5nEkwuojht
PPhmKBYGjwCL1GFJDVPLQtt3ubIkMsy3DeOCOVbBLmxDRMWAnhzTr070hsMzy7AB
uBtF0s85sJRz4wNM1yE+pow1IKYzFM6K1JylsMTeR4lhwvoOQD+bPTUffBA8Vwcx
GpYY31tCtoYK27VfncUrdq//VoHPgDcVg7d4F/obvwQkeEm3tMYxKfNbuuIK0sFx
t/5riYCOMM8pVvxp4Zd78mGnjsyyTmx0DF49yFyAz1bCJcpjgD4zrDwyB0Z9O9nf
fAoJxKhIIhgjrtqG6kg45DF7siiAV3GAZlE7CdIiTag0IcjAhwL9dmV81woCOJP+
oZXbcMk749LJbFX8ANWD98KUgydrEQCFmuzSjluQQDbBRLe9YaRv3cBebgwMH10X
AhHsbJKoCzfArTQLpQL61IrYURt2jothQ3scZswkVVDx6VxzlLlakPEsrPgw2HqZ
KrZIZhLVBRPei1gM0VdzxQYkBr6h9jOFQxIG9oacoccMsp4Hvo/RJ0a7If7YTXty
OEULSWLZ8R+CpUK2imR5THSmu0k5CpBjgNsP6DdpR4KT99CnYZen/bfXDiGOU4xy
lkrXRGVs98LvD8Ee+5FQIKNouyziKiZaQW6ZB1wPM4TLVedz9YT2ONkcMOFkV9Uh
akVmaEBCVN/Ng/BkFjAKWu9zILSgO0FD1mznx6hA2iZwjdRRDYmgZlOvjl/ay8/f
JWDEqxKzQYRFlCaU0IhzKOdbNQs2sFzRtkNriSRyIVyRF8Rt94+z2ntMYHQv4UlM
Nau1ezacsvgZ+X2Yx0KtYKbirFTAJN5whS5Ep1apCQV/o9KsKXjdaWsXXmkOCJrb
S8YZsAMZGBcA9wifbn2cNqtaK0srty5+pRS169GL+0P24/UT/zuQmv8cH+C9UVha
ZKgA49Ms3vUYBObFyalBte3jQHuZ4oA8uwEgP21TW/lG1oD6mnjpLP+UF5thyRzq
mb04MYQQtLF9/45K4+Vv0eycFbGdXAExhqs95BsQTuA9q4YMoYxlUMJ0k6G5ksgA
sxKbsyCqFpncrm/ZakHYRDpZbEDtgDxqH/wv9KKuOKxTpxyRb2CyB+EVVVv8umJA
CvVk1sRI66rcw72blsNYrUO8zsuHe4T3iqlGe8CeVen7RZpJ82enuGEfKcNPzAfe
PB75q3m2q6xKn/DkR4lKMzmvoK4Q0drEnjPVUiFdBOnlKtr8yTEnTk8vhptAEAW7
RhZqVqZ9IY4xNahLlFidICTaYG7O0WeVwvhR76Pv8OcgAybcnyM2+2Z+PbGM5uPx
bzyWS5p48VnV9KydFC9gY0HwXzWsymI8pwoHx7KQuc6gL/tA8E+ptVFnPKew/IsH
KxA5+9r7j4jmPB9pmqO5qy0lNb6iNA0L9VZV0w/51ZBu+mVXWYWEJqou7BE5JU+M
6XGgXEQKorGGxSmou3xBIoROknYN44x4cNwuQ/nrGnzTvSqElSzY4N9sh1wDC7mu
vYMGeAPdhrA20+5bETHAj9q93JGKpK/YlZZQNGsuzwTcpU8wcbA6jS87RP0XOvjR
5Q65xQsX8QITu8LvmiXj5jovXQPUtUdQjJSdPBkDnF3u3pHYtdn8VCgejNcHaKmW
GS1mIulaFCg0gK08O3KFh7KX0slr3IeywzowCarP64Cq5a9ni77O1+wYlM+FazaJ
E/IkGnhmX76dmnOqhHFwSKr+BXtoeVFykscYpj8syYb2pL4eCMyEI+UnugGGT6az
3eVoFfvj+8NB+TIULE7omuknXKnzPDD3LPg1bKeIgLopDaiYfF1rzZORbJ4nBwTr
RvlZHSK7PM3ikZdWQsm4CaqCEki3IOYHjDCBwhrThgKVyDCFdtfk6z8sXFksBBUn
IyXFSVOw/Ps8GEO1D+1/p0nt2UP8hzgPgvjHyLE5sIwzuW+CXNq/cFkw9CbIGGpJ
CWQXhbiYfnRBM773unMG0ZjHsA0jjep5h1xbDefBuHoRcjbAy1HQAN35f+LJyjzV
lnqSxCj21T/Vb9CyS2FIGwuH1glfpPXPalF9qkhRow7ZjHLI2QtUvLKZO+bOcSbL
LroOsKddNd+1O2+UvLz9RadFU1YJNKrk5tGnOuB3T6+0vR8kd+EzxDacFs7nC7u8
VQDLKK4bJprInkIoK6A1d3dU14qfdkJHPEz5q24j/G9GwtYmj6jGxouyUdfkRYqc
ydDjObByRvmkk1AcxXhM6a1z15cX7eUXoCdL4TFM7zctwdIawXefeEUieTrbFmWf
jLA0Y1N8fi1g00ScsG35MRPa8uXl9Q/CGpemX4FqthquVNiPBrs+oaFa81kV0oNv
7JtpgsL8pK74qVtkpDB57GXHd10UR4YOddSOIIR7xt46ZNJHJvOV6LOeFgXHOw2G
no4GtEkSL+0HImy6+G1YKn6n2DQglqzcA7eR4+3tbDn+oR8T6uac7vYWTeYcpSSH
6owXPgzhtK+UQ7Un7d16hYrgS13llXKxzBc+192xiPs/j7FqKlRaUJwHrNz4sKnI
q8YU/wPJHQPGZ1mRomIyUAWLc9pyTgp9Lb00kPLw38kFnb2TPydls064JdrD8d0F
bcFfbElLksQAsSPKpyR6wpFnQrHIG6NTJvl/2Q49fU9fhmnCQ+mwvs1zSxINuVBB
CIuma4LjzyUbR8RIxtEumW5e7W2wyCBl1OmVoZm+WM0k7fiSBHglbkAGarjCo66i
YkZ6ZDoOFe4lXIWJQDJoa/r/rSx3Q0VmL2ktFtZUWp+8ce+gZU4F7VSVQ6piTacP
VcBXTMEf+Pkh46XnfaF1InfeQoksjcTFOe+gH8xER5cxHLTut0B0bo62bREEo0Sa
37K2pHTvBB0OoA7SZjtYhGxYE8f+9+OOCvAG47rhQgT6RPXnUicN3hNB0UDuHsT5
dAscL2em8jE6QsAJIpE1a5pG8kDEv1bCL/LPvDeY2U9S9jy0oGcZFBUnF/0zfTrG
rmZ0FsgK/tKd5FyO9o0S8Gt+e17hv1rQ/eztpG5jC4uYQz8QcfjJPLjrmQqIq8xt
dqI5GUhXv73P56dch0QsNKVYQc8NKpM98qJ46txXY3blE3aWGo+qPALTrtUMiiJ3
tfR8hREUwHiYSBzoBDPvIF3SxjCaC6+0c8C8iKZuocNrc2Tk2TIVxGum6EvHCSuT
IOf/khEcZvOKymi+lX878cwpTPnOPi71OyoiJAW7WY+BuGRdl1UYf/4csNU0Anv0
OsdimWd75do5jqs8+Ir08b6LVuDSicekz4JQCHW293DM+VK3oR4ZLNaPrtHKSiA3
jftOOnCAWRnmMI416dZYzzbNYFKBMP2SKwm80rFJd09bvLiJlRvAcSu8KP5PoPUh
J3ZhfctrDENZLnIa/r+J4tWSOugp7OvoHuekhbX32A7daoORz0TGtPEvpgIPnSNb
zPKrA3ynoqckI1W5ejvOloBTSMBdsB6ld5rrwhQMdnDxUNKuFISR2Th7aJftQR/r
ENHwVX0Gsa8ewlfpLEc7/m7U0Pje95p3RavtCYco+DZ+W87Wbx3ympqVK3Hei8WU
Lo+TfiUEjDJX52/JiiePpfKPDDRxTeivXW4oaHVdRi+BrLAbyNlGy6dPaivihrr6
RxGZ/ACovwcu0ukn7tt1CN0NkmQhheHMAblKHDKmK3q2HKu0008SR13V7dBHl1C+
Iww1BMKrPWXRBqaswJdQAikBf/vOPrNbAZ/2Loc0II4Mhv0YYskhDvk9EKM7oCAt
GoGIUtG3JMTvbMrDWGsNOcAPcA+5nc/mgCFKL3yq5n8F6yYoySNLy8zTgSL8gZ8p
zoNEBk5r5hGPzF8bKFoplP79ts4baLyXoo7pSh26fx+q8L81ijjuheFGNPKfveMc
xHmpYjxf1KLgy0oL7tqJ4QM9G1+YrXcMLrQ1Seg6wthKFTtV/JEQ3m1tcXc03zq4
imWabO+2zUA8AzokhL9fn2RRvFzGzdihthyGqeKy32aTUx6CZ64tGpLFbPHGBboU
6CRS7o1ZY9sH+KSjgJSH+dkJ1vxD0cvZYMaVQWpSnaJSTX1NGQ4VeWWFp82QxxRn
I5/24uPo6hl8+owPm6srzgqQ0eanMMbmBOcjrPHhdMPfziBGDLl/d4HxafROtiVb
i5TGCpWJjy0ls644ec+pOKSxwTZmfLyzqea4FJgQm0vfhdcA0vx5EurmYrxGGxDK
Cze68e82SLTaxHeHjizrHtePrEFCH7/Oj9H0nNN5Wi5caxM4jPcGR98sbQygIWWA
GUVY+2UGyPu4PczDjo02cMKDMqSoEhCEMrGDqhv30JOX7+N+jSOKRU7oPRsnB4ZB
Lwr8hPLpCSJF7nhyqvIf7RXDhQN99o7Zrws3mO+pRUW5B5kSZhnOZHiUDe61lerY
eRByAy9UivGV9ojcN2hWaBpOutMs62o8b0cdN2ySJi5ijqKfnsdM/cseIIb+E8zP
WYAEnLGQlRl3ZKUhpFAOyZDQCtvI3tksQHUBPdKVPLLc5KOHb4tyEZPIVc5DxOIF
nkK6Mt/b/H0oH7MgQHwilVA97kB+GgHlAVZoyT/aiegDq87anetmpm3KezGjX8hw
jfHfNmNEKG4vXHPg7Kcd2OLxPrNtdTcViq8mm3V/mcPTQs//M0L+NCBuGTLtGC6O
0VeZzFLiuUqe5TiD5SKvH/3BFzR3Z3wLJH6DLFWmvh0M9Lb2B23rqKAG+eS0SP8U
VErBzPeeOidp61piLuFbYOPSDiHLmtZKn0ugBckZ3mckBCILF90dtC6dLQxWfJFB
SSJ9mO27C9beEbFZhIP4azxJ8jtkcL6lBcMIT0D9hOvHah18X0dO24z9xu66MORn
ign4bRp6oIk17O3iHIF7DiqIs+7SoByI8Sy6KMl0LYrce1adJSteYlZb95p+Stu9
pF9UJlByPsuikGsxH1Q1avJ3Q9xVVXGR2hMShMyff8B3V8/n0O7aMmC2V5PTuvii
XvZR6Mi1znsRoYGds4/2JbJ7UF6JUlbOejo2m/awWSORhojjHkWxmJSr/jjsymM3
TNudNZv7E67C0cvRSKj1EhkUMkF+6C5OW51+fNuMBFNYfMf9zonLqc5bwf/Rg8ul
4BwvE0iIlAG6rZbESkcYGc8LZoJ+nTSyuALTjV5KYqyhFHLKOjceCcUZpj2qBgnA
+IvXOPzJRnM/kQ2AoGDJzCuvZ4JAmlk/cCSYn1YaiPH8+qTJlQ8xhWm46zC/CHyx
1IiH34zbbAYm+u0Rf4ay+pIb45345JDB469yLy/TAf1K1n6aN0e4q/FPsHtehdyL
q4zSut6WNX7qi93On0dHoJcDzUptEcMbFE0Qd7+R9nt9AL2XiCSv1Y1RJD62JuRd
qP7m91FbTiH0TBac6hnexq/ixRhOm2PN3BBpstyJZixZS5/em3F65aaMyjWS1Bu5
ZJFdiPvd/BCflZKB+fUbfwzwjsHVmlHr3vITZmrL6afy8Qyn2kmEo33Nx0aRZYoI
FKsyCER5AbXWqDPAXUo6Q81nBxFBWnNDXPJOXDCnjBwwnMdOjz2xf+zyl/rQn7wr
iOHF7YA2lnt9VPGftHvVHrrhztWFbLjlZoOT8+xfql/iYjTtBrKi67Vg89zrfgwB
Lch44NqByw1eTql3lbVqHEN6tF1n5QfYMh6X5dPNSikPThUs9r+VGFcW5YEJNUA0
9YXsNaJ+lm0kWqdyN58lCl+V1+5+S8X9MR3qiilWIC8WhaBs6Qfu7saezUlGRA65
EIhEuygSppCqvRLSx5s8FzQXXd8D679iqpJDy4KsEQfSYT6hQ03xVBhYyCT6qRZf
p54/6BezGFQyUOLqQi5nQEF3o3oHPIHmlOkPTZLHaxzLIDyy6hnQw4K5GEwuOSqn
zPV1blXaGdpvH0l2ejHGjzZuwb/WIrbrMeHd+Is1WTQTRqoPMZR68F0fdrXegZxt
763UA4gxLy+vUGeHacQsE3MMTXD6Y6cR1ISQwNbmvt3r1aqgLnQKt86ir1ZGjS9x
UongTCbmT3hm+Ga9tvIro4OBTvC7ELyDKnceFW1Rp6i6TJP/u5lULmqYZpUsDGbu
ryFSEIcK1StEmhUbCerwwHy2JGG3Ema8gxcvoiR+KYQNcdIvt5046PKyEgOv2c5i
fB0PFnnCD/p+QsGRDczz9jWCeRRWWv9sD2gjwUx9prKrxQHiEr65Bcd0RQOmj9bM
tTc+zGmzQaQZtDCoYwCO5sMrQvMsAYeDAZvjNtzKdmaDZK9bdlJhJmdvzVIjkr/E
BEKt0m0Iqt/CtWjOacOjjP01MVKUCnUEA2KLo8DQsO9njjHbROoHcfkr3VprMGm+
BEBySAahBWxPQrpsgGIikGanwtQmtF3+9sXtzoUvkTQ/2/RtOnZzU8hUzkSs4OoR
7O/NMdXGjwHAl2L8DQh5J1CivPP5JLmgmxI0v090lzL2GXcwVTM+5UPlY1ZlnlSO
xQWpVN6VkVpE+APxeWW2PhudwRtlP23isYToriNxNEvRbf8rjIxLtPnZ24P6IEWC
Ut4Vm3j2YppCj1GS3OPVLBJWb+2JrG2eEJPTp8bgT/f5KcpsRA0gKqWm7Hi4+mYH
qOFNiuG3yYplZUXwA/pzo+62Q+WPBMjOZ2c0+UyhInklI6mCyQW3lK9RSZZnQ+9P
Rcc06tpQvnf0CsraOGJjqd606ownyLo6wpbnzMKhnMKf+Ht1/e1240jn8hXM9aI9
9A5dqgdJzJq8UaRyx+WOhB+OZN/u8YIKVw14RdbP5nC0QEDdU7KCCovkGAoOj1Bz
L3w/bEaXHBEFMVa6vC/e5XfZo3UPoJ9X+/KTCJGkH194asbOlR6mX8rH/uZvf3oR
txLySiFpaLYS2Pfe7qcR65sbL7ZUArDo5AjxNo4dvenLg99GdywnyIk5uYgeNrcd
sChC/S1wkOdVzJ1XooKUrMgwq40eoZvYUazkSuEUclslaIrVOYl6c9m2RxPIvPvN
3n+OyHSNjHF0A2fspTSCrgCPsEYAIgf/z25VnCNDE/mzD06hTs1eTJs4LUPGrc4E
eNDdUdAYAVf4FqQIkGApvjtiELJqU9BOhqWlzJKRfI/qtcas1ifuTvthNvCwdPFq
Yt+WEHv0fKpiZ99N7gxq0jTv7cXo7jaA/BNF4tIneO68Gtctv6uXVzZTG58jUp44
fSVTYp7I8vM8Ww82aYuo+2s4P4zjEXmBBuvQKKCf4/XPp3QeGuEaCVSBOd1/9+QE
WsCSyh/nSHlJkFKzxcmDpseGgNUzTSuu7YcYTwum5F+QvFIC66P/YDTy3xdkh1T3
7e8L5gjHzf3kqmvgwkHtnv+7/x75ltVFsMWnC91rbcfbf/V8hWHVPppoNoktOMnC
Sd1oStOvrxsf91ApGOO2oIoIQoHiRAPWetedcKV3CuJy04eVbYOflMg7IXMa3W8I
TeF/uH0uOQ/aBkm5i3WBbnYFjKgPR8Rbqcfvb0NUqWFdxY2m9G6tU0nw5qb6nrI5
9JroF3+1ohkZ5S/bzh6dVTEWMol88IC+6fKhp9k7I7u4DhAbpPknhGEdtxHqwmhX
n3ZGUJ2qb7B10lU0OBsG7vsbOSVtBwAygQkQVl02+8NP4jkmM0pnBr14+ztxR5rQ
lBvuPzGeAQxIuMQOpmkcKEV+AQV9fO9m+HHk2Q3RwuYjdKzeUxRwPj23SiLJZM/y
ypvejVpspR4zN09qN+2mvyc5nUX+adLnXd2db5NX8EbBfJUNTmsSXTQoK5YlxKf4
w5OvyvrRoaRMzlXVW0uGpnMxSNYDw0rP4T1BqwGyXXeAAWch5Kh9gYNWjOVCmVdt
la4xTv96qHX3hYZEutfBpDbtBUqaEJq4C7u1JWaoVl8SHPxumV5kdDnjFd+06alr
G07yaJi95VxiGx4hqMDUt+DuIRaFCFv4SyeBeqaJIZc9i7kFsihv+n+qhAmyRvGF
8vdaJcKaDS3MiRPv+ncdppdIiBdp/a5XwNkUBpx/Om/KH5ACC+e/T2V1ysV9GX/P
YHYU4gpK6zYfdcQ3RWOJnM4le/YP43eeDi65ahxGU6Zalmty5L/mrFsMedAUs8in
xwDU8fsnzGT0Up9jDc+XgK2E3B2X7xhLPx5jGY7rgnJ/JI9v+S94mowIzF8NjikR
I9w4nXcuVsOTbU4EcSfRgJb3xEGLiWO1yqCnySaSIDPBXDf1ei9USm03ljBDuu/m
df8vh9WnS0zuF/DLDM/NV1edeesLXN/pm4UdgsbGVA8/rnDcoI98IFrrdCm610Ou
4KJar8fMzU+43Eu2JossgpUprLXBrNFilYiiBgcoB+wc+yfnHP7ub/oLz4kmSKSk
aW8JPHtOqbKOfAqUHCFf1J3X2cznEExuIq5PiYw2AJviWuG0Hwp5GbfPZqhuAD85
grE9VuasuIRilT8NEG7Eful33UX/qskckfwHHQ8lSzKFB22B3SweiUafL3sX2C84
oprhHgxToFTJ8Akq7+5wUVMzQH2W9Pv/1jRNIIxWr/Je0QEoQaFcacr/tspaY19x
OOs6NzugrFAoGJ9uD5gRPf2Wy6Az6Qve51iLkaCl+TKECPcicwBHzh2sKie0v0OI
nwcfeNjci75nUo5BX7JKDfNQT6fKgX6DLslEBwHYD9xNA9mIal1TnVBUU0gsWB4X
G8FdvvqBSYvHA9Lj/lrh28O8faGpXa8YLmuexHRd47QnV9ppN/Rbbv+15YF9lqju
/W0txrG/67uiXt+O++kw9MbV5oD3tr2G2yi31IWGJMqtTO5obZpJYlgG7MxsQ2G3
QmwVJFHtRTZ+kAxZg6GS7GN6P7l/HSEG2uLqNfhSgJntABTDobRlqEuisbCRray4
qgakE73CmSEPewI0tKqMcXAAEeRokr3Sj1k/VDUA1k2VrP6gRZdwpX1fvgOAroVr
pS57aO22Mg4W4cM//XzYjU9uHNmTKWiHLaMMBoyHnVD3FZsfgztOrxn8swQuFTHu
7BIJ+zdrYyhzF116kvZ0Bs+NuA8hdBbySxeU5NPBIaXUbSBZ+OkJeElKeFANR6FC
zBy1Dvu5GXecivzc27LOYBmWfhfQj7LS0DslObLIydyl08MmH2sXr4IkHWDKtsml
72e+8XjmQGcN56hDDYS9vdenXL5c1A/fALZmEmvHNfp33Tm5anirOjgg3Gukduem
BXSuWREVF6Sj1r+sFAy/BkiaXk5dsf2Q31HqYd3/F4jY7z8etgy8HzvLtEqUrUu3
PPLhJRTFSpAS/0J7bJ5gSG1Z6ofHHiqFuJr9kJKRK8NCxcewPazxuIa+1ygb7L8r
D4x5OaZhsVnTEWQ4OTh9vE6AsHowEGE6bRJXvhVltlrbAZLpag+FpQETMkpFMpEw
m+kuVD8VuJ1xl/MmU8NwWV65rVfUYNsrrfb5RLd24tlBjccvvjD+y+mOKM8Gh58q
LAkZQfST59pKcXv2S9SrfgjIGH0aW8ywZT60EAKF6oDqErNmTtK3C35uonXFbgU3
iBZDneLFkfw4rIgIW4wt6AeKewkMjrOc09UnQKQsRx61NTFqw6l1FIcBYpMnczCi
gqvSJztLpDTYSHSPkTlNnL1CPyM63f/f6qRXVB8Mfnh0e+C7BPu3vx9Xy9eLGz0F
VOobZJWsMkrfKRpXEC+Yn7iPFyOL1TdjZB3wlTnXLsdkWiIkIQVtWiTya8RUn7AG
tMUlUdj5yDFk4eqz3VbWABpbbGwWgwHsu67vQT2Jqr1+xfQA5nPi+gP5uzXKGCze
9csou5NANdyM0mTYZMLmpmTyQbieh16Oqje6Ax05w9kRaVihXomPHskaL83ckBqk
zIzQSzV+o38iHVyIFWsdUdTADOOXetR8/cjLu6033DNOOOEhxNVVfW2Wd89C2Opx
IGGj2vE3Fom2bzua0hWhRjeQcTJSCuSYqn0JI3gi1wyT5E4GAuhriQdLwULqJ++j
zxoXqzj65kRuaNB3/fCI1vXHX/9aFz3iHCux+2lxsSlNPR6OZWmPVIUxugKfbPj4
6Fh54xN6CMRBhiZQz1Qc41xeuJ7sY9maqOeuO+OWHQO90syLiMqAAbGcFkOfRcqD
77XNHYP84KnpMcw5g/6aw35fbABeT/UoqYTcFs6du6AGBjAProkZyFdU7fvw+Hsp
sN9CBNy7xvHY7SZfAgObj/EvYUjd2GFJGsU3naERbc3TiL4A3hNhFyLOgD1XeHrM
nzRC+Np6HAuR0c8Hu2kTgBnE7A9G/yxZK1d3C0GZZLylNYKj8p1N41jKi4A4W805
asCVSSU7CijbirnrDHGoIdLOHAbk4wbhe/lCTFZ0Gzh6Y+Tv/rYHWESPxPKVA3s6
pk4Y9yc4yq706YV+REwvBpgnZ1aMHix4MLuZHF0B2wosU7H5qoGPiu0LwiHNAKr4
9ViPUz5XkL5eG84ywEnQ6mMWc0ebPGNk1vMKlddUFwzOitemvNlpeRvUkpd5ZBvp
sesQjVlO8PoIeTpqNeOp7OIHu26Bt8utdMJDBhhY/w+5tZ2OaZ6nBluEYb3hc8LY
G7B/k1DHgAMG/JydAfrZkm6p5NsHSCJtfcDBQgwhFT2HhB5xjQUD7iEBldpijN5D
NZ/ZH5UUTp0J0dJtAsP6KreVxbUrFBQtN6DxOkMr60XGC5a09ScDtojzQ3OX+XVN
GSV0E+3KLbRIpDLRNORIOTV6+Wk6ksRXtnh7ekY/1FUdTx9s68RE5cOP6Jl52im+
xYpT0ZhEjDqVTb0FcLLlnuWXaWTAI7IQOvfezxgvIFIs3LHQHDpRwI30dYxT7uyz
Hi8LrLwsg5JzpZf79UqMKaulguo0LIINinold2J076pX+nxnGQXRfMegvPjYnNmT
FnK9FZk1bPbHAX7RSiIJjx0N+3OR246uVB5u3M9AbO+sdSjCRfr3NDlgD97F7b2B
jsJrXLjW0BYiSTQQjKW6IoCVtIoN0kZ8Mgnld9wKBEcQhaSzkZBiC/olluGh+w/R
Ub1g7185g98FCw+/Z0skyjt9nMxtyPkzrWC8QJC51mP5VpGBC40bCCLO7galn6fC
`pragma protect end_protected

endmodule
